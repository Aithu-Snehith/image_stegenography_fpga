module	helloworld(i_clk,
			o_ledg,
			i_rts, i_uart_rx, o_cts,
			o_uart_tx);
	//
	input		i_clk;
	output	wire	o_ledg;
	input		i_rts, i_uart_rx;
	output		o_cts;
	output	wire	o_uart_tx;

	assign	o_cts = 1'b1;

	// If i_setup isnt set up as an input parameter, it needs to be set.
	// We do so here, to a setting appropriate to create a 115200 Baud
	// comms system from a 100MHz clock.  This also sets us to an 8-bit
	// data word, 1-stop bit, and no parity.
	wire	[29:0]	i_setup;
	assign		i_setup = 30'd868;	// 115200 Baud, if clk @ 100MHz

	reg	pwr_reset;
	initial	pwr_reset = 1'b1;
	always @(posedge i_clk)
		pwr_reset <= 1'b0;

	reg	[24:0]	ledctr;
	initial	ledctr = 0;
	always @(posedge i_clk)
		if (!o_uart_tx)
			ledctr <= 0;
		else if (ledctr != {(25){1'b1}})
			ledctr <= ledctr + 1'b1;
	assign	o_ledg = !ledctr[24];

 reg[119:0] message;
 	initial message = 120'b011100110110111001100101011010000110100101110100011010000010000001101001011100110010000001101000011001010111001001100101;

	reg [7:0] img [0:4095]

	initial begin
		img[4095] = 8'b00011000;
		img[4094] = 8'b00010110;
		img[4093] = 8'b10100000;
		img[4092] = 8'b01111111;
		img[4091] = 8'b11001010;
		img[4090] = 8'b11100101;
		img[4089] = 8'b11111000;
		img[4088] = 8'b10101011;
		img[4087] = 8'b10110010;
		img[4086] = 8'b11010100;
		img[4085] = 8'b11001110;
		img[4084] = 8'b11001000;
		img[4083] = 8'b10011111;
		img[4082] = 8'b10000000;
		img[4081] = 8'b10001011;
		img[4080] = 8'b10011100;
		img[4079] = 8'b10101010;
		img[4078] = 8'b10111011;
		img[4077] = 8'b10100100;
		img[4076] = 8'b01100010;
		img[4075] = 8'b00011101;
		img[4074] = 8'b00000000;
		img[4073] = 8'b00011010;
		img[4072] = 8'b00100000;
		img[4071] = 8'b01001011;
		img[4070] = 8'b00000000;
		img[4069] = 8'b00000000;
		img[4068] = 8'b00001011;
		img[4067] = 8'b00000000;
		img[4066] = 8'b00010100;
		img[4065] = 8'b00000011;
		img[4064] = 8'b00010000;
		img[4063] = 8'b00000110;
		img[4062] = 8'b00001110;
		img[4061] = 8'b00000000;
		img[4060] = 8'b00000010;
		img[4059] = 8'b00000110;
		img[4058] = 8'b00000110;
		img[4057] = 8'b00010010;
		img[4056] = 8'b00010011;
		img[4055] = 8'b00100100;
		img[4054] = 8'b00010100;
		img[4053] = 8'b00001111;
		img[4052] = 8'b00010001;
		img[4051] = 8'b00010000;
		img[4050] = 8'b00010100;
		img[4049] = 8'b00010110;
		img[4048] = 8'b00010101;
		img[4047] = 8'b00100101;
		img[4046] = 8'b00011010;
		img[4045] = 8'b00001110;
		img[4044] = 8'b00010110;
		img[4043] = 8'b00010011;
		img[4042] = 8'b00010000;
		img[4041] = 8'b00010101;
		img[4040] = 8'b00010101;
		img[4039] = 8'b00000100;
		img[4038] = 8'b00010011;
		img[4037] = 8'b00000110;
		img[4036] = 8'b00000110;
		img[4035] = 8'b00000000;
		img[4034] = 8'b00011000;
		img[4033] = 8'b00101001;
		img[4032] = 8'b00000100;
		img[4031] = 8'b10000100;
		img[4030] = 8'b11000110;
		img[4029] = 8'b10011001;
		img[4028] = 8'b00111100;
		img[4027] = 8'b01101000;
		img[4026] = 8'b01100100;
		img[4025] = 8'b01110010;
		img[4024] = 8'b10001000;
		img[4023] = 8'b10111101;
		img[4022] = 8'b11101101;
		img[4021] = 8'b01101000;
		img[4020] = 8'b10001001;
		img[4019] = 8'b10001101;
		img[4018] = 8'b10100010;
		img[4017] = 8'b01111101;
		img[4016] = 8'b01100100;
		img[4015] = 8'b01101001;
		img[4014] = 8'b01101000;
		img[4013] = 8'b10000011;
		img[4012] = 8'b01010110;
		img[4011] = 8'b00111110;
		img[4010] = 8'b00101101;
		img[4009] = 8'b00011010;
		img[4008] = 8'b00111111;
		img[4007] = 8'b00011111;
		img[4006] = 8'b00011000;
		img[4005] = 8'b00000000;
		img[4004] = 8'b00000011;
		img[4003] = 8'b00000010;
		img[4002] = 8'b00011101;
		img[4001] = 8'b00101011;
		img[4000] = 8'b00000001;
		img[3999] = 8'b00001011;
		img[3998] = 8'b00010100;
		img[3997] = 8'b00001011;
		img[3996] = 8'b00001000;
		img[3995] = 8'b00000101;
		img[3994] = 8'b00010011;
		img[3993] = 8'b00010111;
		img[3992] = 8'b00011001;
		img[3991] = 8'b00001111;
		img[3990] = 8'b00011110;
		img[3989] = 8'b00000111;
		img[3988] = 8'b00001010;
		img[3987] = 8'b00011101;
		img[3986] = 8'b00010010;
		img[3985] = 8'b00010001;
		img[3984] = 8'b00010010;
		img[3983] = 8'b00010110;
		img[3982] = 8'b00101111;
		img[3981] = 8'b00000000;
		img[3980] = 8'b00010011;
		img[3979] = 8'b00001101;
		img[3978] = 8'b00011010;
		img[3977] = 8'b00010110;
		img[3976] = 8'b00011001;
		img[3975] = 8'b00001101;
		img[3974] = 8'b00000010;
		img[3973] = 8'b00001001;
		img[3972] = 8'b00000101;
		img[3971] = 8'b00000101;
		img[3970] = 8'b00011001;
		img[3969] = 8'b00001100;
		img[3968] = 8'b00010100;
		img[3967] = 8'b01100111;
		img[3966] = 8'b01110111;
		img[3965] = 8'b00010110;
		img[3964] = 8'b01110110;
		img[3963] = 8'b01110101;
		img[3962] = 8'b01101101;
		img[3961] = 8'b01010101;
		img[3960] = 8'b10000011;
		img[3959] = 8'b11000111;
		img[3958] = 8'b10000010;
		img[3957] = 8'b01001110;
		img[3956] = 8'b00111101;
		img[3955] = 8'b01011111;
		img[3954] = 8'b01101000;
		img[3953] = 8'b01100101;
		img[3952] = 8'b01000111;
		img[3951] = 8'b01010011;
		img[3950] = 8'b01101000;
		img[3949] = 8'b01111010;
		img[3948] = 8'b01111001;
		img[3947] = 8'b00111000;
		img[3946] = 8'b00101100;
		img[3945] = 8'b00100100;
		img[3944] = 8'b01100000;
		img[3943] = 8'b00110001;
		img[3942] = 8'b00000000;
		img[3941] = 8'b00000100;
		img[3940] = 8'b00001010;
		img[3939] = 8'b00011110;
		img[3938] = 8'b00010110;
		img[3937] = 8'b00011001;
		img[3936] = 8'b00010101;
		img[3935] = 8'b00100111;
		img[3934] = 8'b00000011;
		img[3933] = 8'b00001111;
		img[3932] = 8'b00011011;
		img[3931] = 8'b00010011;
		img[3930] = 8'b00100101;
		img[3929] = 8'b00000000;
		img[3928] = 8'b00110001;
		img[3927] = 8'b00000001;
		img[3926] = 8'b00011000;
		img[3925] = 8'b00000000;
		img[3924] = 8'b00000010;
		img[3923] = 8'b00010111;
		img[3922] = 8'b00100001;
		img[3921] = 8'b00001110;
		img[3920] = 8'b00011110;
		img[3919] = 8'b00011110;
		img[3918] = 8'b00000000;
		img[3917] = 8'b00001111;
		img[3916] = 8'b00010100;
		img[3915] = 8'b00010101;
		img[3914] = 8'b00000000;
		img[3913] = 8'b00011101;
		img[3912] = 8'b00011000;
		img[3911] = 8'b00010100;
		img[3910] = 8'b00100000;
		img[3909] = 8'b00000000;
		img[3908] = 8'b00010001;
		img[3907] = 8'b00001011;
		img[3906] = 8'b00010100;
		img[3905] = 8'b00100001;
		img[3904] = 8'b00000100;
		img[3903] = 8'b01001111;
		img[3902] = 8'b01010000;
		img[3901] = 8'b01011110;
		img[3900] = 8'b01100000;
		img[3899] = 8'b01101101;
		img[3898] = 8'b01111001;
		img[3897] = 8'b01111111;
		img[3896] = 8'b10001011;
		img[3895] = 8'b10010001;
		img[3894] = 8'b01000101;
		img[3893] = 8'b01000111;
		img[3892] = 8'b01010101;
		img[3891] = 8'b01010111;
		img[3890] = 8'b01101110;
		img[3889] = 8'b01010001;
		img[3888] = 8'b01010100;
		img[3887] = 8'b01101001;
		img[3886] = 8'b01101110;
		img[3885] = 8'b01111001;
		img[3884] = 8'b01100001;
		img[3883] = 8'b01000100;
		img[3882] = 8'b00101011;
		img[3881] = 8'b00111001;
		img[3880] = 8'b01110110;
		img[3879] = 8'b00111000;
		img[3878] = 8'b00010001;
		img[3877] = 8'b00101010;
		img[3876] = 8'b00101010;
		img[3875] = 8'b00011000;
		img[3874] = 8'b00001011;
		img[3873] = 8'b00110000;
		img[3872] = 8'b00001110;
		img[3871] = 8'b00010000;
		img[3870] = 8'b00010010;
		img[3869] = 8'b00101011;
		img[3868] = 8'b01000010;
		img[3867] = 8'b00001101;
		img[3866] = 8'b00101000;
		img[3865] = 8'b00110100;
		img[3864] = 8'b00010011;
		img[3863] = 8'b00000000;
		img[3862] = 8'b00000000;
		img[3861] = 8'b00000101;
		img[3860] = 8'b00000000;
		img[3859] = 8'b00000000;
		img[3858] = 8'b00010111;
		img[3857] = 8'b00010110;
		img[3856] = 8'b00001000;
		img[3855] = 8'b00001101;
		img[3854] = 8'b00001010;
		img[3853] = 8'b00010110;
		img[3852] = 8'b00011010;
		img[3851] = 8'b00000000;
		img[3850] = 8'b00010000;
		img[3849] = 8'b00010001;
		img[3848] = 8'b00001110;
		img[3847] = 8'b00100001;
		img[3846] = 8'b00000010;
		img[3845] = 8'b00001000;
		img[3844] = 8'b00000001;
		img[3843] = 8'b00000000;
		img[3842] = 8'b00000110;
		img[3841] = 8'b00000000;
		img[3840] = 8'b00000001;
		img[3839] = 8'b01000100;
		img[3838] = 8'b00001010;
		img[3837] = 8'b00010001;
		img[3836] = 8'b00100100;
		img[3835] = 8'b00100110;
		img[3834] = 8'b00101101;
		img[3833] = 8'b00110000;
		img[3832] = 8'b01001010;
		img[3831] = 8'b01111001;
		img[3830] = 8'b01000000;
		img[3829] = 8'b01000101;
		img[3828] = 8'b00111001;
		img[3827] = 8'b01001100;
		img[3826] = 8'b01101110;
		img[3825] = 8'b01110001;
		img[3824] = 8'b01001011;
		img[3823] = 8'b01011010;
		img[3822] = 8'b01100110;
		img[3821] = 8'b01101000;
		img[3820] = 8'b01111000;
		img[3819] = 8'b01000100;
		img[3818] = 8'b01000011;
		img[3817] = 8'b01111110;
		img[3816] = 8'b01010110;
		img[3815] = 8'b01010000;
		img[3814] = 8'b00111111;
		img[3813] = 8'b00100111;
		img[3812] = 8'b00101000;
		img[3811] = 8'b00010001;
		img[3810] = 8'b00011110;
		img[3809] = 8'b00101000;
		img[3808] = 8'b00011100;
		img[3807] = 8'b00101100;
		img[3806] = 8'b00100110;
		img[3805] = 8'b00010010;
		img[3804] = 8'b00111101;
		img[3803] = 8'b01010000;
		img[3802] = 8'b01100111;
		img[3801] = 8'b00101110;
		img[3800] = 8'b00011011;
		img[3799] = 8'b00001010;
		img[3798] = 8'b00001111;
		img[3797] = 8'b00001000;
		img[3796] = 8'b00010011;
		img[3795] = 8'b00010101;
		img[3794] = 8'b00001000;
		img[3793] = 8'b00100011;
		img[3792] = 8'b00000110;
		img[3791] = 8'b00011001;
		img[3790] = 8'b00001101;
		img[3789] = 8'b00000111;
		img[3788] = 8'b00011101;
		img[3787] = 8'b00000111;
		img[3786] = 8'b00010000;
		img[3785] = 8'b00101000;
		img[3784] = 8'b00000001;
		img[3783] = 8'b00011011;
		img[3782] = 8'b00001111;
		img[3781] = 8'b00000110;
		img[3780] = 8'b00000000;
		img[3779] = 8'b00000111;
		img[3778] = 8'b00000111;
		img[3777] = 8'b00000000;
		img[3776] = 8'b00000010;
		img[3775] = 8'b01011001;
		img[3774] = 8'b00100101;
		img[3773] = 8'b00111111;
		img[3772] = 8'b00011010;
		img[3771] = 8'b00000010;
		img[3770] = 8'b00000000;
		img[3769] = 8'b00000000;
		img[3768] = 8'b00000000;
		img[3767] = 8'b00000001;
		img[3766] = 8'b00011001;
		img[3765] = 8'b00100000;
		img[3764] = 8'b00110000;
		img[3763] = 8'b00110111;
		img[3762] = 8'b01001110;
		img[3761] = 8'b01011011;
		img[3760] = 8'b01001000;
		img[3759] = 8'b01000011;
		img[3758] = 8'b01011001;
		img[3757] = 8'b01010101;
		img[3756] = 8'b01011101;
		img[3755] = 8'b00100100;
		img[3754] = 8'b01011010;
		img[3753] = 8'b01100011;
		img[3752] = 8'b01101010;
		img[3751] = 8'b01110000;
		img[3750] = 8'b01010010;
		img[3749] = 8'b00000100;
		img[3748] = 8'b00000111;
		img[3747] = 8'b00001011;
		img[3746] = 8'b00101110;
		img[3745] = 8'b00100111;
		img[3744] = 8'b00011111;
		img[3743] = 8'b00101101;
		img[3742] = 8'b00101100;
		img[3741] = 8'b01001010;
		img[3740] = 8'b10001010;
		img[3739] = 8'b01001001;
		img[3738] = 8'b00111111;
		img[3737] = 8'b01101001;
		img[3736] = 8'b00011011;
		img[3735] = 8'b00101010;
		img[3734] = 8'b00010010;
		img[3733] = 8'b00010111;
		img[3732] = 8'b00001001;
		img[3731] = 8'b00000100;
		img[3730] = 8'b00000101;
		img[3729] = 8'b00000110;
		img[3728] = 8'b00010101;
		img[3727] = 8'b00010000;
		img[3726] = 8'b00001011;
		img[3725] = 8'b00010010;
		img[3724] = 8'b00011011;
		img[3723] = 8'b00000000;
		img[3722] = 8'b00011001;
		img[3721] = 8'b00001000;
		img[3720] = 8'b00010001;
		img[3719] = 8'b00000000;
		img[3718] = 8'b00000000;
		img[3717] = 8'b00001000;
		img[3716] = 8'b00000000;
		img[3715] = 8'b00001000;
		img[3714] = 8'b00011111;
		img[3713] = 8'b00001011;
		img[3712] = 8'b00001011;
		img[3711] = 8'b01001111;
		img[3710] = 8'b01000001;
		img[3709] = 8'b00110100;
		img[3708] = 8'b00101011;
		img[3707] = 8'b00000111;
		img[3706] = 8'b00001101;
		img[3705] = 8'b00010101;
		img[3704] = 8'b00000001;
		img[3703] = 8'b00000000;
		img[3702] = 8'b00000000;
		img[3701] = 8'b00000011;
		img[3700] = 8'b00000001;
		img[3699] = 8'b00010001;
		img[3698] = 8'b00101000;
		img[3697] = 8'b00101011;
		img[3696] = 8'b01000100;
		img[3695] = 8'b01001101;
		img[3694] = 8'b01111110;
		img[3693] = 8'b01100100;
		img[3692] = 8'b01001001;
		img[3691] = 8'b01011101;
		img[3690] = 8'b01101000;
		img[3689] = 8'b01100111;
		img[3688] = 8'b01100110;
		img[3687] = 8'b01001110;
		img[3686] = 8'b01001011;
		img[3685] = 8'b00011111;
		img[3684] = 8'b00000110;
		img[3683] = 8'b00001010;
		img[3682] = 8'b00011011;
		img[3681] = 8'b00100100;
		img[3680] = 8'b01000111;
		img[3679] = 8'b01011000;
		img[3678] = 8'b00011010;
		img[3677] = 8'b00110111;
		img[3676] = 8'b01010101;
		img[3675] = 8'b00101010;
		img[3674] = 8'b01110000;
		img[3673] = 8'b01011110;
		img[3672] = 8'b01000010;
		img[3671] = 8'b00100010;
		img[3670] = 8'b00101001;
		img[3669] = 8'b00111010;
		img[3668] = 8'b00011011;
		img[3667] = 8'b00100111;
		img[3666] = 8'b00011010;
		img[3665] = 8'b00001000;
		img[3664] = 8'b00100010;
		img[3663] = 8'b00010100;
		img[3662] = 8'b00001110;
		img[3661] = 8'b00000110;
		img[3660] = 8'b00000110;
		img[3659] = 8'b00001110;
		img[3658] = 8'b00001001;
		img[3657] = 8'b00000000;
		img[3656] = 8'b00000010;
		img[3655] = 8'b00000000;
		img[3654] = 8'b00001011;
		img[3653] = 8'b00000110;
		img[3652] = 8'b00000000;
		img[3651] = 8'b00011101;
		img[3650] = 8'b00000000;
		img[3649] = 8'b00000011;
		img[3648] = 8'b00011000;
		img[3647] = 8'b01101101;
		img[3646] = 8'b00011001;
		img[3645] = 8'b01101010;
		img[3644] = 8'b00100111;
		img[3643] = 8'b00010101;
		img[3642] = 8'b00000110;
		img[3641] = 8'b00000111;
		img[3640] = 8'b00010111;
		img[3639] = 8'b00001001;
		img[3638] = 8'b00000000;
		img[3637] = 8'b00010100;
		img[3636] = 8'b00000000;
		img[3635] = 8'b00000000;
		img[3634] = 8'b00000000;
		img[3633] = 8'b00000101;
		img[3632] = 8'b00000111;
		img[3631] = 8'b01011011;
		img[3630] = 8'b01001011;
		img[3629] = 8'b00100111;
		img[3628] = 8'b00101100;
		img[3627] = 8'b01000101;
		img[3626] = 8'b00111111;
		img[3625] = 8'b01011011;
		img[3624] = 8'b10000101;
		img[3623] = 8'b01010010;
		img[3622] = 8'b00101101;
		img[3621] = 8'b00011111;
		img[3620] = 8'b00010111;
		img[3619] = 8'b00011110;
		img[3618] = 8'b00110001;
		img[3617] = 8'b01000110;
		img[3616] = 8'b01011000;
		img[3615] = 8'b01001100;
		img[3614] = 8'b01010011;
		img[3613] = 8'b01011110;
		img[3612] = 8'b01000110;
		img[3611] = 8'b01011110;
		img[3610] = 8'b01111000;
		img[3609] = 8'b01111111;
		img[3608] = 8'b01010000;
		img[3607] = 8'b01001111;
		img[3606] = 8'b01001000;
		img[3605] = 8'b00100111;
		img[3604] = 8'b00110100;
		img[3603] = 8'b00101101;
		img[3602] = 8'b00001011;
		img[3601] = 8'b00000100;
		img[3600] = 8'b00001100;
		img[3599] = 8'b00001111;
		img[3598] = 8'b00000111;
		img[3597] = 8'b00000100;
		img[3596] = 8'b00000000;
		img[3595] = 8'b00000000;
		img[3594] = 8'b00001001;
		img[3593] = 8'b00000111;
		img[3592] = 8'b00001011;
		img[3591] = 8'b00000000;
		img[3590] = 8'b00010110;
		img[3589] = 8'b00001001;
		img[3588] = 8'b00011011;
		img[3587] = 8'b00000000;
		img[3586] = 8'b00000000;
		img[3585] = 8'b00001100;
		img[3584] = 8'b00001111;
		img[3583] = 8'b01010110;
		img[3582] = 8'b01110110;
		img[3581] = 8'b10001011;
		img[3580] = 8'b01000001;
		img[3579] = 8'b00100000;
		img[3578] = 8'b00010000;
		img[3577] = 8'b00011011;
		img[3576] = 8'b00001011;
		img[3575] = 8'b00001101;
		img[3574] = 8'b00000000;
		img[3573] = 8'b00000000;
		img[3572] = 8'b00010011;
		img[3571] = 8'b00001100;
		img[3570] = 8'b00001011;
		img[3569] = 8'b00000011;
		img[3568] = 8'b00000001;
		img[3567] = 8'b00000000;
		img[3566] = 8'b00000100;
		img[3565] = 8'b00100010;
		img[3564] = 8'b00110011;
		img[3563] = 8'b00110101;
		img[3562] = 8'b00111111;
		img[3561] = 8'b01011010;
		img[3560] = 8'b10000010;
		img[3559] = 8'b10001001;
		img[3558] = 8'b01011101;
		img[3557] = 8'b00111111;
		img[3556] = 8'b00011101;
		img[3555] = 8'b01000000;
		img[3554] = 8'b00110000;
		img[3553] = 8'b01010001;
		img[3552] = 8'b01010110;
		img[3551] = 8'b10000010;
		img[3550] = 8'b01101001;
		img[3549] = 8'b10001100;
		img[3548] = 8'b01100010;
		img[3547] = 8'b01111100;
		img[3546] = 8'b01101111;
		img[3545] = 8'b10001110;
		img[3544] = 8'b10011110;
		img[3543] = 8'b01010011;
		img[3542] = 8'b01101101;
		img[3541] = 8'b00101100;
		img[3540] = 8'b00110101;
		img[3539] = 8'b00110100;
		img[3538] = 8'b00010101;
		img[3537] = 8'b00001101;
		img[3536] = 8'b00000000;
		img[3535] = 8'b00011011;
		img[3534] = 8'b00000000;
		img[3533] = 8'b00001010;
		img[3532] = 8'b00001001;
		img[3531] = 8'b00000010;
		img[3530] = 8'b00001011;
		img[3529] = 8'b00001001;
		img[3528] = 8'b00100010;
		img[3527] = 8'b00000100;
		img[3526] = 8'b00001100;
		img[3525] = 8'b00000000;
		img[3524] = 8'b00001000;
		img[3523] = 8'b00001101;
		img[3522] = 8'b00001101;
		img[3521] = 8'b00001100;
		img[3520] = 8'b00010000;
		img[3519] = 8'b10111101;
		img[3518] = 8'b10111011;
		img[3517] = 8'b10001010;
		img[3516] = 8'b01000110;
		img[3515] = 8'b01000101;
		img[3514] = 8'b00100010;
		img[3513] = 8'b00000111;
		img[3512] = 8'b00001010;
		img[3511] = 8'b00000001;
		img[3510] = 8'b00000000;
		img[3509] = 8'b00001011;
		img[3508] = 8'b00010100;
		img[3507] = 8'b00000110;
		img[3506] = 8'b00001110;
		img[3505] = 8'b00001010;
		img[3504] = 8'b00011010;
		img[3503] = 8'b00000000;
		img[3502] = 8'b00000000;
		img[3501] = 8'b00000000;
		img[3500] = 8'b00000011;
		img[3499] = 8'b01001001;
		img[3498] = 8'b00101111;
		img[3497] = 8'b01101110;
		img[3496] = 8'b10001001;
		img[3495] = 8'b10001000;
		img[3494] = 8'b01001001;
		img[3493] = 8'b10000110;
		img[3492] = 8'b00110101;
		img[3491] = 8'b01001010;
		img[3490] = 8'b01101111;
		img[3489] = 8'b01001001;
		img[3488] = 8'b01100001;
		img[3487] = 8'b10001000;
		img[3486] = 8'b10000110;
		img[3485] = 8'b10000001;
		img[3484] = 8'b10010011;
		img[3483] = 8'b10010000;
		img[3482] = 8'b10001001;
		img[3481] = 8'b10010101;
		img[3480] = 8'b10011000;
		img[3479] = 8'b01110100;
		img[3478] = 8'b01100111;
		img[3477] = 8'b01110100;
		img[3476] = 8'b01100001;
		img[3475] = 8'b00101110;
		img[3474] = 8'b00011000;
		img[3473] = 8'b00000000;
		img[3472] = 8'b00010111;
		img[3471] = 8'b00001111;
		img[3470] = 8'b00000110;
		img[3469] = 8'b00010011;
		img[3468] = 8'b00000000;
		img[3467] = 8'b00010001;
		img[3466] = 8'b00000011;
		img[3465] = 8'b00000001;
		img[3464] = 8'b00010011;
		img[3463] = 8'b00000111;
		img[3462] = 8'b00011010;
		img[3461] = 8'b00001001;
		img[3460] = 8'b00001011;
		img[3459] = 8'b00000001;
		img[3458] = 8'b00100100;
		img[3457] = 8'b00000011;
		img[3456] = 8'b00000000;
		img[3455] = 8'b00011011;
		img[3454] = 8'b01011101;
		img[3453] = 8'b10001001;
		img[3452] = 8'b01111000;
		img[3451] = 8'b01100011;
		img[3450] = 8'b00011011;
		img[3449] = 8'b00000011;
		img[3448] = 8'b00001111;
		img[3447] = 8'b00001101;
		img[3446] = 8'b00000000;
		img[3445] = 8'b00010110;
		img[3444] = 8'b00000000;
		img[3443] = 8'b00000000;
		img[3442] = 8'b00000000;
		img[3441] = 8'b00000000;
		img[3440] = 8'b00001001;
		img[3439] = 8'b00010000;
		img[3438] = 8'b00000000;
		img[3437] = 8'b00000000;
		img[3436] = 8'b00001001;
		img[3435] = 8'b00000010;
		img[3434] = 8'b00111011;
		img[3433] = 8'b01011111;
		img[3432] = 8'b00111001;
		img[3431] = 8'b01101000;
		img[3430] = 8'b01110000;
		img[3429] = 8'b01001111;
		img[3428] = 8'b01001111;
		img[3427] = 8'b10000100;
		img[3426] = 8'b01100011;
		img[3425] = 8'b01010011;
		img[3424] = 8'b01110110;
		img[3423] = 8'b01111100;
		img[3422] = 8'b01111000;
		img[3421] = 8'b10100100;
		img[3420] = 8'b10010000;
		img[3419] = 8'b10011100;
		img[3418] = 8'b10011100;
		img[3417] = 8'b10010000;
		img[3416] = 8'b10010010;
		img[3415] = 8'b01101000;
		img[3414] = 8'b01110110;
		img[3413] = 8'b01110001;
		img[3412] = 8'b01011000;
		img[3411] = 8'b00110111;
		img[3410] = 8'b00100001;
		img[3409] = 8'b00100011;
		img[3408] = 8'b00101010;
		img[3407] = 8'b00100001;
		img[3406] = 8'b00001011;
		img[3405] = 8'b00100110;
		img[3404] = 8'b00011001;
		img[3403] = 8'b00010000;
		img[3402] = 8'b00001000;
		img[3401] = 8'b00000000;
		img[3400] = 8'b00010101;
		img[3399] = 8'b00010101;
		img[3398] = 8'b00010001;
		img[3397] = 8'b00011001;
		img[3396] = 8'b00000000;
		img[3395] = 8'b00010011;
		img[3394] = 8'b00000000;
		img[3393] = 8'b00001011;
		img[3392] = 8'b00000000;
		img[3391] = 8'b10001010;
		img[3390] = 8'b10010010;
		img[3389] = 8'b10000100;
		img[3388] = 8'b10001101;
		img[3387] = 8'b01111010;
		img[3386] = 8'b01010000;
		img[3385] = 8'b01100011;
		img[3384] = 8'b00011110;
		img[3383] = 8'b00001100;
		img[3382] = 8'b00000000;
		img[3381] = 8'b00001110;
		img[3380] = 8'b00010100;
		img[3379] = 8'b00001010;
		img[3378] = 8'b00000000;
		img[3377] = 8'b00001011;
		img[3376] = 8'b00000110;
		img[3375] = 8'b00001011;
		img[3374] = 8'b00000010;
		img[3373] = 8'b00000000;
		img[3372] = 8'b00001001;
		img[3371] = 8'b00000000;
		img[3370] = 8'b00001010;
		img[3369] = 8'b00011111;
		img[3368] = 8'b01011010;
		img[3367] = 8'b10100001;
		img[3366] = 8'b10001000;
		img[3365] = 8'b01111001;
		img[3364] = 8'b10010110;
		img[3363] = 8'b10100001;
		img[3362] = 8'b10010011;
		img[3361] = 8'b01100101;
		img[3360] = 8'b10001110;
		img[3359] = 8'b10001010;
		img[3358] = 8'b10010000;
		img[3357] = 8'b10001110;
		img[3356] = 8'b10010110;
		img[3355] = 8'b10010000;
		img[3354] = 8'b10010110;
		img[3353] = 8'b10011000;
		img[3352] = 8'b10011100;
		img[3351] = 8'b10010110;
		img[3350] = 8'b10000000;
		img[3349] = 8'b10000111;
		img[3348] = 8'b01100011;
		img[3347] = 8'b01000011;
		img[3346] = 8'b01010001;
		img[3345] = 8'b00100111;
		img[3344] = 8'b00110100;
		img[3343] = 8'b00101110;
		img[3342] = 8'b00010001;
		img[3341] = 8'b00111011;
		img[3340] = 8'b00010111;
		img[3339] = 8'b00001100;
		img[3338] = 8'b00000100;
		img[3337] = 8'b00001100;
		img[3336] = 8'b00001000;
		img[3335] = 8'b00010110;
		img[3334] = 8'b00000001;
		img[3333] = 8'b00000000;
		img[3332] = 8'b00010101;
		img[3331] = 8'b00001101;
		img[3330] = 8'b00011101;
		img[3329] = 8'b00000000;
		img[3328] = 8'b00000011;
		img[3327] = 8'b10111010;
		img[3326] = 8'b10000110;
		img[3325] = 8'b10011000;
		img[3324] = 8'b10011100;
		img[3323] = 8'b10000011;
		img[3322] = 8'b10010100;
		img[3321] = 8'b01111110;
		img[3320] = 8'b01010011;
		img[3319] = 8'b00100110;
		img[3318] = 8'b00001110;
		img[3317] = 8'b00010000;
		img[3316] = 8'b00000000;
		img[3315] = 8'b00001110;
		img[3314] = 8'b00001101;
		img[3313] = 8'b00010101;
		img[3312] = 8'b00000000;
		img[3311] = 8'b00011000;
		img[3310] = 8'b00000000;
		img[3309] = 8'b00000110;
		img[3308] = 8'b00001001;
		img[3307] = 8'b00010111;
		img[3306] = 8'b00000101;
		img[3305] = 8'b00101101;
		img[3304] = 8'b01011111;
		img[3303] = 8'b10000000;
		img[3302] = 8'b10011100;
		img[3301] = 8'b10011010;
		img[3300] = 8'b10011101;
		img[3299] = 8'b10010111;
		img[3298] = 8'b10011111;
		img[3297] = 8'b10011111;
		img[3296] = 8'b10010111;
		img[3295] = 8'b01111011;
		img[3294] = 8'b10001110;
		img[3293] = 8'b10001000;
		img[3292] = 8'b10011000;
		img[3291] = 8'b10010011;
		img[3290] = 8'b10010001;
		img[3289] = 8'b10010101;
		img[3288] = 8'b10010000;
		img[3287] = 8'b10001111;
		img[3286] = 8'b10011000;
		img[3285] = 8'b10010100;
		img[3284] = 8'b10010111;
		img[3283] = 8'b01101000;
		img[3282] = 8'b01011010;
		img[3281] = 8'b00101100;
		img[3280] = 8'b01000101;
		img[3279] = 8'b00110011;
		img[3278] = 8'b00110011;
		img[3277] = 8'b01000010;
		img[3276] = 8'b00011101;
		img[3275] = 8'b00100000;
		img[3274] = 8'b00000011;
		img[3273] = 8'b00010001;
		img[3272] = 8'b00000000;
		img[3271] = 8'b00000100;
		img[3270] = 8'b00000001;
		img[3269] = 8'b00010011;
		img[3268] = 8'b00001001;
		img[3267] = 8'b00000010;
		img[3266] = 8'b00010010;
		img[3265] = 8'b00001100;
		img[3264] = 8'b00000000;
		img[3263] = 8'b10001010;
		img[3262] = 8'b10001000;
		img[3261] = 8'b10100010;
		img[3260] = 8'b11000100;
		img[3259] = 8'b10111110;
		img[3258] = 8'b10010010;
		img[3257] = 8'b01101000;
		img[3256] = 8'b00111101;
		img[3255] = 8'b00011000;
		img[3254] = 8'b00001010;
		img[3253] = 8'b00001000;
		img[3252] = 8'b00000111;
		img[3251] = 8'b00010011;
		img[3250] = 8'b00000110;
		img[3249] = 8'b00000011;
		img[3248] = 8'b00000111;
		img[3247] = 8'b00000100;
		img[3246] = 8'b00000000;
		img[3245] = 8'b00000000;
		img[3244] = 8'b00001111;
		img[3243] = 8'b00000011;
		img[3242] = 8'b00100110;
		img[3241] = 8'b00111110;
		img[3240] = 8'b01010111;
		img[3239] = 8'b00110110;
		img[3238] = 8'b10011100;
		img[3237] = 8'b10010110;
		img[3236] = 8'b10010110;
		img[3235] = 8'b10010000;
		img[3234] = 8'b10010110;
		img[3233] = 8'b10010011;
		img[3232] = 8'b10010001;
		img[3231] = 8'b01101111;
		img[3230] = 8'b10001100;
		img[3229] = 8'b10000011;
		img[3228] = 8'b10010001;
		img[3227] = 8'b10001000;
		img[3226] = 8'b10010100;
		img[3225] = 8'b10010111;
		img[3224] = 8'b10010010;
		img[3223] = 8'b10010011;
		img[3222] = 8'b10001110;
		img[3221] = 8'b10001011;
		img[3220] = 8'b10001110;
		img[3219] = 8'b10011001;
		img[3218] = 8'b01001111;
		img[3217] = 8'b01110111;
		img[3216] = 8'b01101111;
		img[3215] = 8'b00110011;
		img[3214] = 8'b01100101;
		img[3213] = 8'b00101100;
		img[3212] = 8'b00101010;
		img[3211] = 8'b00101001;
		img[3210] = 8'b00000000;
		img[3209] = 8'b00010101;
		img[3208] = 8'b00001110;
		img[3207] = 8'b00010101;
		img[3206] = 8'b00001000;
		img[3205] = 8'b00000000;
		img[3204] = 8'b00001010;
		img[3203] = 8'b00000011;
		img[3202] = 8'b00000110;
		img[3201] = 8'b00001010;
		img[3200] = 8'b00001000;
		img[3199] = 8'b10110010;
		img[3198] = 8'b10101000;
		img[3197] = 8'b10111010;
		img[3196] = 8'b10000100;
		img[3195] = 8'b11011010;
		img[3194] = 8'b10011001;
		img[3193] = 8'b10010110;
		img[3192] = 8'b00110110;
		img[3191] = 8'b00011111;
		img[3190] = 8'b00011110;
		img[3189] = 8'b00000001;
		img[3188] = 8'b00001011;
		img[3187] = 8'b00001101;
		img[3186] = 8'b00000111;
		img[3185] = 8'b00010000;
		img[3184] = 8'b00000000;
		img[3183] = 8'b00010001;
		img[3182] = 8'b00001001;
		img[3181] = 8'b00000000;
		img[3180] = 8'b00001000;
		img[3179] = 8'b00011100;
		img[3178] = 8'b00000110;
		img[3177] = 8'b01101000;
		img[3176] = 8'b01010010;
		img[3175] = 8'b10010010;
		img[3174] = 8'b10011010;
		img[3173] = 8'b10010111;
		img[3172] = 8'b10001011;
		img[3171] = 8'b10100000;
		img[3170] = 8'b10011000;
		img[3169] = 8'b10011011;
		img[3168] = 8'b01111000;
		img[3167] = 8'b10010101;
		img[3166] = 8'b10011000;
		img[3165] = 8'b10010010;
		img[3164] = 8'b10010101;
		img[3163] = 8'b10010010;
		img[3162] = 8'b10001110;
		img[3161] = 8'b10000111;
		img[3160] = 8'b10000110;
		img[3159] = 8'b10001110;
		img[3158] = 8'b10001101;
		img[3157] = 8'b10000110;
		img[3156] = 8'b10001111;
		img[3155] = 8'b10010011;
		img[3154] = 8'b01010101;
		img[3153] = 8'b01111000;
		img[3152] = 8'b10001100;
		img[3151] = 8'b01100010;
		img[3150] = 8'b01100110;
		img[3149] = 8'b01010111;
		img[3148] = 8'b00111110;
		img[3147] = 8'b00011100;
		img[3146] = 8'b00001011;
		img[3145] = 8'b00100001;
		img[3144] = 8'b00001100;
		img[3143] = 8'b00010000;
		img[3142] = 8'b00001001;
		img[3141] = 8'b00000000;
		img[3140] = 8'b00000101;
		img[3139] = 8'b00001110;
		img[3138] = 8'b00011001;
		img[3137] = 8'b00010001;
		img[3136] = 8'b00010011;
		img[3135] = 8'b00010100;
		img[3134] = 8'b00101001;
		img[3133] = 8'b00100111;
		img[3132] = 8'b01011001;
		img[3131] = 8'b01100111;
		img[3130] = 8'b00111001;
		img[3129] = 8'b01110001;
		img[3128] = 8'b01101101;
		img[3127] = 8'b01100001;
		img[3126] = 8'b00011110;
		img[3125] = 8'b00001000;
		img[3124] = 8'b00010000;
		img[3123] = 8'b00001101;
		img[3122] = 8'b00001111;
		img[3121] = 8'b00001110;
		img[3120] = 8'b00010010;
		img[3119] = 8'b00011000;
		img[3118] = 8'b00000001;
		img[3117] = 8'b00001111;
		img[3116] = 8'b00010000;
		img[3115] = 8'b00101001;
		img[3114] = 8'b00100101;
		img[3113] = 8'b00011001;
		img[3112] = 8'b01100001;
		img[3111] = 8'b10010111;
		img[3110] = 8'b10010100;
		img[3109] = 8'b01111110;
		img[3108] = 8'b01110000;
		img[3107] = 8'b01110111;
		img[3106] = 8'b10000111;
		img[3105] = 8'b10010100;
		img[3104] = 8'b10010000;
		img[3103] = 8'b01110111;
		img[3102] = 8'b10001001;
		img[3101] = 8'b10010100;
		img[3100] = 8'b10010001;
		img[3099] = 8'b10010110;
		img[3098] = 8'b10010100;
		img[3097] = 8'b10010111;
		img[3096] = 8'b10010110;
		img[3095] = 8'b10010001;
		img[3094] = 8'b10000111;
		img[3093] = 8'b10000010;
		img[3092] = 8'b01111100;
		img[3091] = 8'b01100110;
		img[3090] = 8'b01101010;
		img[3089] = 8'b10001110;
		img[3088] = 8'b10000011;
		img[3087] = 8'b01000111;
		img[3086] = 8'b01011111;
		img[3085] = 8'b01010000;
		img[3084] = 8'b01010001;
		img[3083] = 8'b01011000;
		img[3082] = 8'b00101010;
		img[3081] = 8'b00110010;
		img[3080] = 8'b00011001;
		img[3079] = 8'b00000111;
		img[3078] = 8'b00001111;
		img[3077] = 8'b00000000;
		img[3076] = 8'b00000010;
		img[3075] = 8'b00100000;
		img[3074] = 8'b00001010;
		img[3073] = 8'b00010010;
		img[3072] = 8'b00010011;
		img[3071] = 8'b00001001;
		img[3070] = 8'b00000000;
		img[3069] = 8'b00001010;
		img[3068] = 8'b00000000;
		img[3067] = 8'b00100011;
		img[3066] = 8'b00111110;
		img[3065] = 8'b01010101;
		img[3064] = 8'b01001100;
		img[3063] = 8'b01001000;
		img[3062] = 8'b00011110;
		img[3061] = 8'b00010000;
		img[3060] = 8'b00011100;
		img[3059] = 8'b00001100;
		img[3058] = 8'b00000000;
		img[3057] = 8'b00001011;
		img[3056] = 8'b00000111;
		img[3055] = 8'b00010111;
		img[3054] = 8'b00001110;
		img[3053] = 8'b01011010;
		img[3052] = 8'b00100000;
		img[3051] = 8'b00100010;
		img[3050] = 8'b00001010;
		img[3049] = 8'b00101000;
		img[3048] = 8'b01000001;
		img[3047] = 8'b01101101;
		img[3046] = 8'b10010010;
		img[3045] = 8'b10101010;
		img[3044] = 8'b10101001;
		img[3043] = 8'b10001101;
		img[3042] = 8'b01111111;
		img[3041] = 8'b01111011;
		img[3040] = 8'b10010101;
		img[3039] = 8'b10001011;
		img[3038] = 8'b10010001;
		img[3037] = 8'b10001001;
		img[3036] = 8'b10000011;
		img[3035] = 8'b10001110;
		img[3034] = 8'b10001011;
		img[3033] = 8'b10000010;
		img[3032] = 8'b10000101;
		img[3031] = 8'b10001100;
		img[3030] = 8'b10000101;
		img[3029] = 8'b01111111;
		img[3028] = 8'b10000000;
		img[3027] = 8'b01101011;
		img[3026] = 8'b10001001;
		img[3025] = 8'b10000010;
		img[3024] = 8'b10000001;
		img[3023] = 8'b10001110;
		img[3022] = 8'b01110001;
		img[3021] = 8'b01010110;
		img[3020] = 8'b01111111;
		img[3019] = 8'b01111010;
		img[3018] = 8'b10000010;
		img[3017] = 8'b01010110;
		img[3016] = 8'b01001001;
		img[3015] = 8'b00001110;
		img[3014] = 8'b00010000;
		img[3013] = 8'b00010010;
		img[3012] = 8'b00100010;
		img[3011] = 8'b00001001;
		img[3010] = 8'b00000111;
		img[3009] = 8'b00010100;
		img[3008] = 8'b00001100;
		img[3007] = 8'b00011000;
		img[3006] = 8'b00010110;
		img[3005] = 8'b00001101;
		img[3004] = 8'b00001011;
		img[3003] = 8'b00000000;
		img[3002] = 8'b00000010;
		img[3001] = 8'b00011000;
		img[3000] = 8'b00101101;
		img[2999] = 8'b01110010;
		img[2998] = 8'b01011100;
		img[2997] = 8'b01000001;
		img[2996] = 8'b00011101;
		img[2995] = 8'b00010111;
		img[2994] = 8'b00001100;
		img[2993] = 8'b00010100;
		img[2992] = 8'b00001111;
		img[2991] = 8'b00000100;
		img[2990] = 8'b00001101;
		img[2989] = 8'b01000010;
		img[2988] = 8'b00011110;
		img[2987] = 8'b00011110;
		img[2986] = 8'b00010110;
		img[2985] = 8'b00110101;
		img[2984] = 8'b00110001;
		img[2983] = 8'b01001000;
		img[2982] = 8'b01001000;
		img[2981] = 8'b01001011;
		img[2980] = 8'b01011000;
		img[2979] = 8'b01101011;
		img[2978] = 8'b01111110;
		img[2977] = 8'b10010011;
		img[2976] = 8'b10011110;
		img[2975] = 8'b10110100;
		img[2974] = 8'b10111000;
		img[2973] = 8'b10001000;
		img[2972] = 8'b10001011;
		img[2971] = 8'b10001111;
		img[2970] = 8'b10001101;
		img[2969] = 8'b10001110;
		img[2968] = 8'b10001001;
		img[2967] = 8'b10001000;
		img[2966] = 8'b10010011;
		img[2965] = 8'b10001011;
		img[2964] = 8'b10001011;
		img[2963] = 8'b10001110;
		img[2962] = 8'b10000011;
		img[2961] = 8'b01111100;
		img[2960] = 8'b10000011;
		img[2959] = 8'b10001001;
		img[2958] = 8'b10000100;
		img[2957] = 8'b01100100;
		img[2956] = 8'b01111110;
		img[2955] = 8'b10010000;
		img[2954] = 8'b10100101;
		img[2953] = 8'b10000011;
		img[2952] = 8'b01010000;
		img[2951] = 8'b00000000;
		img[2950] = 8'b00001000;
		img[2949] = 8'b00000000;
		img[2948] = 8'b00011011;
		img[2947] = 8'b00000101;
		img[2946] = 8'b00010011;
		img[2945] = 8'b00010110;
		img[2944] = 8'b00000001;
		img[2943] = 8'b00101101;
		img[2942] = 8'b00011001;
		img[2941] = 8'b00010110;
		img[2940] = 8'b00011010;
		img[2939] = 8'b00100011;
		img[2938] = 8'b00101011;
		img[2937] = 8'b00010111;
		img[2936] = 8'b00001111;
		img[2935] = 8'b00010100;
		img[2934] = 8'b01001001;
		img[2933] = 8'b01000010;
		img[2932] = 8'b00111000;
		img[2931] = 8'b00100011;
		img[2930] = 8'b00101110;
		img[2929] = 8'b00100011;
		img[2928] = 8'b00100101;
		img[2927] = 8'b00000000;
		img[2926] = 8'b00001100;
		img[2925] = 8'b00011010;
		img[2924] = 8'b00010010;
		img[2923] = 8'b00000101;
		img[2922] = 8'b00001111;
		img[2921] = 8'b00010100;
		img[2920] = 8'b00011001;
		img[2919] = 8'b00100001;
		img[2918] = 8'b00010110;
		img[2917] = 8'b00001101;
		img[2916] = 8'b00001010;
		img[2915] = 8'b00010100;
		img[2914] = 8'b00101110;
		img[2913] = 8'b01000111;
		img[2912] = 8'b01101010;
		img[2911] = 8'b01111011;
		img[2910] = 8'b01110001;
		img[2909] = 8'b10000001;
		img[2908] = 8'b10001100;
		img[2907] = 8'b10001001;
		img[2906] = 8'b10010101;
		img[2905] = 8'b10001101;
		img[2904] = 8'b10001100;
		img[2903] = 8'b10010000;
		img[2902] = 8'b10001000;
		img[2901] = 8'b01111000;
		img[2900] = 8'b01111001;
		img[2899] = 8'b10000101;
		img[2898] = 8'b10010000;
		img[2897] = 8'b10011111;
		img[2896] = 8'b10010101;
		img[2895] = 8'b10100101;
		img[2894] = 8'b10100111;
		img[2893] = 8'b10001010;
		img[2892] = 8'b01110001;
		img[2891] = 8'b01111000;
		img[2890] = 8'b01011111;
		img[2889] = 8'b10001001;
		img[2888] = 8'b00111001;
		img[2887] = 8'b00000100;
		img[2886] = 8'b00000000;
		img[2885] = 8'b00000001;
		img[2884] = 8'b00010001;
		img[2883] = 8'b00001100;
		img[2882] = 8'b00000010;
		img[2881] = 8'b00000000;
		img[2880] = 8'b00001111;
		img[2879] = 8'b00010100;
		img[2878] = 8'b00010111;
		img[2877] = 8'b00010100;
		img[2876] = 8'b00001000;
		img[2875] = 8'b00001001;
		img[2874] = 8'b00001011;
		img[2873] = 8'b00100001;
		img[2872] = 8'b00011101;
		img[2871] = 8'b00001011;
		img[2870] = 8'b00000000;
		img[2869] = 8'b00101001;
		img[2868] = 8'b00100001;
		img[2867] = 8'b00010000;
		img[2866] = 8'b00101110;
		img[2865] = 8'b00110111;
		img[2864] = 8'b00010101;
		img[2863] = 8'b00000101;
		img[2862] = 8'b00010010;
		img[2861] = 8'b00010111;
		img[2860] = 8'b00011011;
		img[2859] = 8'b00001011;
		img[2858] = 8'b00100100;
		img[2857] = 8'b00000000;
		img[2856] = 8'b00010001;
		img[2855] = 8'b00000001;
		img[2854] = 8'b00010010;
		img[2853] = 8'b00000111;
		img[2852] = 8'b00000000;
		img[2851] = 8'b00000000;
		img[2850] = 8'b00000011;
		img[2849] = 8'b00000000;
		img[2848] = 8'b00010110;
		img[2847] = 8'b01010011;
		img[2846] = 8'b10000110;
		img[2845] = 8'b10011011;
		img[2844] = 8'b10011010;
		img[2843] = 8'b10100011;
		img[2842] = 8'b10011000;
		img[2841] = 8'b10101110;
		img[2840] = 8'b10111101;
		img[2839] = 8'b11000000;
		img[2838] = 8'b10100111;
		img[2837] = 8'b10101000;
		img[2836] = 8'b10011001;
		img[2835] = 8'b10100011;
		img[2834] = 8'b01011000;
		img[2833] = 8'b00100010;
		img[2832] = 8'b01100010;
		img[2831] = 8'b10001001;
		img[2830] = 8'b10000000;
		img[2829] = 8'b01111100;
		img[2828] = 8'b10111000;
		img[2827] = 8'b11000000;
		img[2826] = 8'b10011110;
		img[2825] = 8'b01011111;
		img[2824] = 8'b01001100;
		img[2823] = 8'b00101100;
		img[2822] = 8'b00000000;
		img[2821] = 8'b00000000;
		img[2820] = 8'b00101011;
		img[2819] = 8'b00000000;
		img[2818] = 8'b00001100;
		img[2817] = 8'b00000000;
		img[2816] = 8'b00011011;
		img[2815] = 8'b00010100;
		img[2814] = 8'b00100010;
		img[2813] = 8'b00010010;
		img[2812] = 8'b00011110;
		img[2811] = 8'b00000011;
		img[2810] = 8'b00001101;
		img[2809] = 8'b00001010;
		img[2808] = 8'b00000110;
		img[2807] = 8'b00010000;
		img[2806] = 8'b00100001;
		img[2805] = 8'b00001010;
		img[2804] = 8'b00010010;
		img[2803] = 8'b00000111;
		img[2802] = 8'b00001100;
		img[2801] = 8'b00111101;
		img[2800] = 8'b00010100;
		img[2799] = 8'b01010011;
		img[2798] = 8'b00110111;
		img[2797] = 8'b00000000;
		img[2796] = 8'b00000100;
		img[2795] = 8'b00000000;
		img[2794] = 8'b00000010;
		img[2793] = 8'b00000000;
		img[2792] = 8'b00000000;
		img[2791] = 8'b00010000;
		img[2790] = 8'b00001010;
		img[2789] = 8'b00000100;
		img[2788] = 8'b00000000;
		img[2787] = 8'b00000000;
		img[2786] = 8'b00000110;
		img[2785] = 8'b00000000;
		img[2784] = 8'b00011000;
		img[2783] = 8'b00010100;
		img[2782] = 8'b01111100;
		img[2781] = 8'b10010110;
		img[2780] = 8'b11010011;
		img[2779] = 8'b10101001;
		img[2778] = 8'b11000000;
		img[2777] = 8'b11000000;
		img[2776] = 8'b10100011;
		img[2775] = 8'b10010100;
		img[2774] = 8'b10000001;
		img[2773] = 8'b10000010;
		img[2772] = 8'b10110010;
		img[2771] = 8'b10001111;
		img[2770] = 8'b10001011;
		img[2769] = 8'b10000000;
		img[2768] = 8'b10100001;
		img[2767] = 8'b01110111;
		img[2766] = 8'b01101001;
		img[2765] = 8'b01000001;
		img[2764] = 8'b10010101;
		img[2763] = 8'b01111001;
		img[2762] = 8'b10110110;
		img[2761] = 8'b01101110;
		img[2760] = 8'b00011011;
		img[2759] = 8'b00101110;
		img[2758] = 8'b00001010;
		img[2757] = 8'b00000000;
		img[2756] = 8'b00001000;
		img[2755] = 8'b00001000;
		img[2754] = 8'b00000000;
		img[2753] = 8'b00000000;
		img[2752] = 8'b00000010;
		img[2751] = 8'b00001010;
		img[2750] = 8'b00010001;
		img[2749] = 8'b00100000;
		img[2748] = 8'b00011010;
		img[2747] = 8'b00001111;
		img[2746] = 8'b00001010;
		img[2745] = 8'b00000100;
		img[2744] = 8'b00000001;
		img[2743] = 8'b00010000;
		img[2742] = 8'b00001010;
		img[2741] = 8'b00110011;
		img[2740] = 8'b01000000;
		img[2739] = 8'b00101110;
		img[2738] = 8'b00110011;
		img[2737] = 8'b01100001;
		img[2736] = 8'b01000101;
		img[2735] = 8'b01001111;
		img[2734] = 8'b01010100;
		img[2733] = 8'b01001100;
		img[2732] = 8'b00011000;
		img[2731] = 8'b00011000;
		img[2730] = 8'b00010111;
		img[2729] = 8'b00011100;
		img[2728] = 8'b00001001;
		img[2727] = 8'b00000000;
		img[2726] = 8'b00000011;
		img[2725] = 8'b00000000;
		img[2724] = 8'b00000000;
		img[2723] = 8'b00010101;
		img[2722] = 8'b00000110;
		img[2721] = 8'b00100000;
		img[2720] = 8'b00010011;
		img[2719] = 8'b00001010;
		img[2718] = 8'b01010000;
		img[2717] = 8'b00111000;
		img[2716] = 8'b01011001;
		img[2715] = 8'b01110100;
		img[2714] = 8'b01101110;
		img[2713] = 8'b01101010;
		img[2712] = 8'b10100101;
		img[2711] = 8'b10010000;
		img[2710] = 8'b10010001;
		img[2709] = 8'b11010001;
		img[2708] = 8'b10011101;
		img[2707] = 8'b10100011;
		img[2706] = 8'b10100001;
		img[2705] = 8'b10011000;
		img[2704] = 8'b10001011;
		img[2703] = 8'b00100010;
		img[2702] = 8'b00111101;
		img[2701] = 8'b01001011;
		img[2700] = 8'b01010011;
		img[2699] = 8'b00111101;
		img[2698] = 8'b01010100;
		img[2697] = 8'b01111010;
		img[2696] = 8'b00101010;
		img[2695] = 8'b00001101;
		img[2694] = 8'b00000000;
		img[2693] = 8'b00001100;
		img[2692] = 8'b00010010;
		img[2691] = 8'b00000101;
		img[2690] = 8'b00001011;
		img[2689] = 8'b00000110;
		img[2688] = 8'b00000110;
		img[2687] = 8'b00010110;
		img[2686] = 8'b00001111;
		img[2685] = 8'b00000000;
		img[2684] = 8'b00001001;
		img[2683] = 8'b00001011;
		img[2682] = 8'b00010110;
		img[2681] = 8'b00011010;
		img[2680] = 8'b00010001;
		img[2679] = 8'b00011101;
		img[2678] = 8'b00000000;
		img[2677] = 8'b00000010;
		img[2676] = 8'b00010100;
		img[2675] = 8'b00101111;
		img[2674] = 8'b00101001;
		img[2673] = 8'b01001000;
		img[2672] = 8'b01000100;
		img[2671] = 8'b00110010;
		img[2670] = 8'b00110010;
		img[2669] = 8'b00010100;
		img[2668] = 8'b00010000;
		img[2667] = 8'b00100100;
		img[2666] = 8'b00001110;
		img[2665] = 8'b00010110;
		img[2664] = 8'b00000000;
		img[2663] = 8'b00010011;
		img[2662] = 8'b00011011;
		img[2661] = 8'b00000000;
		img[2660] = 8'b00010000;
		img[2659] = 8'b00010111;
		img[2658] = 8'b00101010;
		img[2657] = 8'b00100101;
		img[2656] = 8'b00000111;
		img[2655] = 8'b00011010;
		img[2654] = 8'b00000000;
		img[2653] = 8'b00010001;
		img[2652] = 8'b00100100;
		img[2651] = 8'b00110111;
		img[2650] = 8'b01011101;
		img[2649] = 8'b01100010;
		img[2648] = 8'b01111100;
		img[2647] = 8'b01110111;
		img[2646] = 8'b01110010;
		img[2645] = 8'b10110001;
		img[2644] = 8'b10011000;
		img[2643] = 8'b11000101;
		img[2642] = 8'b10000111;
		img[2641] = 8'b10110100;
		img[2640] = 8'b10001111;
		img[2639] = 8'b00001001;
		img[2638] = 8'b00000000;
		img[2637] = 8'b00110000;
		img[2636] = 8'b00000001;
		img[2635] = 8'b00001111;
		img[2634] = 8'b00001010;
		img[2633] = 8'b00110001;
		img[2632] = 8'b00110011;
		img[2631] = 8'b00001001;
		img[2630] = 8'b00001010;
		img[2629] = 8'b00011000;
		img[2628] = 8'b00001000;
		img[2627] = 8'b00000011;
		img[2626] = 8'b00001111;
		img[2625] = 8'b00010010;
		img[2624] = 8'b00000000;
		img[2623] = 8'b00101110;
		img[2622] = 8'b00001001;
		img[2621] = 8'b00000000;
		img[2620] = 8'b00000000;
		img[2619] = 8'b00010011;
		img[2618] = 8'b00010101;
		img[2617] = 8'b00010100;
		img[2616] = 8'b00010010;
		img[2615] = 8'b00000111;
		img[2614] = 8'b00000011;
		img[2613] = 8'b00011000;
		img[2612] = 8'b00000110;
		img[2611] = 8'b00000011;
		img[2610] = 8'b00000100;
		img[2609] = 8'b00001101;
		img[2608] = 8'b00000011;
		img[2607] = 8'b00000101;
		img[2606] = 8'b00000101;
		img[2605] = 8'b00101100;
		img[2604] = 8'b00100011;
		img[2603] = 8'b00000011;
		img[2602] = 8'b00010010;
		img[2601] = 8'b00000010;
		img[2600] = 8'b00010111;
		img[2599] = 8'b00000100;
		img[2598] = 8'b00000000;
		img[2597] = 8'b00011000;
		img[2596] = 8'b00010011;
		img[2595] = 8'b00100011;
		img[2594] = 8'b00010111;
		img[2593] = 8'b00001100;
		img[2592] = 8'b00010010;
		img[2591] = 8'b00100010;
		img[2590] = 8'b00000010;
		img[2589] = 8'b00000000;
		img[2588] = 8'b00001110;
		img[2587] = 8'b00000010;
		img[2586] = 8'b00001101;
		img[2585] = 8'b00110111;
		img[2584] = 8'b01010111;
		img[2583] = 8'b10010110;
		img[2582] = 8'b10000101;
		img[2581] = 8'b10100010;
		img[2580] = 8'b10010110;
		img[2579] = 8'b10001000;
		img[2578] = 8'b10011111;
		img[2577] = 8'b10100010;
		img[2576] = 8'b10001000;
		img[2575] = 8'b00010011;
		img[2574] = 8'b00011000;
		img[2573] = 8'b00010010;
		img[2572] = 8'b00001100;
		img[2571] = 8'b00011001;
		img[2570] = 8'b00110010;
		img[2569] = 8'b01010101;
		img[2568] = 8'b01010001;
		img[2567] = 8'b00000100;
		img[2566] = 8'b00000000;
		img[2565] = 8'b00000010;
		img[2564] = 8'b00000000;
		img[2563] = 8'b00000000;
		img[2562] = 8'b00000111;
		img[2561] = 8'b00000000;
		img[2560] = 8'b00000000;
		img[2559] = 8'b00011011;
		img[2558] = 8'b00010000;
		img[2557] = 8'b00000101;
		img[2556] = 8'b00001111;
		img[2555] = 8'b00100011;
		img[2554] = 8'b00000000;
		img[2553] = 8'b00001011;
		img[2552] = 8'b00001000;
		img[2551] = 8'b00001100;
		img[2550] = 8'b00001110;
		img[2549] = 8'b00001010;
		img[2548] = 8'b00010111;
		img[2547] = 8'b00010111;
		img[2546] = 8'b00000000;
		img[2545] = 8'b00000000;
		img[2544] = 8'b00000000;
		img[2543] = 8'b00000111;
		img[2542] = 8'b00000000;
		img[2541] = 8'b00001111;
		img[2540] = 8'b00011011;
		img[2539] = 8'b00000000;
		img[2538] = 8'b00000011;
		img[2537] = 8'b00001011;
		img[2536] = 8'b00001000;
		img[2535] = 8'b00000000;
		img[2534] = 8'b00000010;
		img[2533] = 8'b00000010;
		img[2532] = 8'b00000011;
		img[2531] = 8'b00000000;
		img[2530] = 8'b00011010;
		img[2529] = 8'b00000000;
		img[2528] = 8'b00011011;
		img[2527] = 8'b00011111;
		img[2526] = 8'b00001011;
		img[2525] = 8'b00000111;
		img[2524] = 8'b00010010;
		img[2523] = 8'b00001111;
		img[2522] = 8'b00001000;
		img[2521] = 8'b00000010;
		img[2520] = 8'b00000001;
		img[2519] = 8'b00011111;
		img[2518] = 8'b01000000;
		img[2517] = 8'b01011011;
		img[2516] = 8'b01111111;
		img[2515] = 8'b10010100;
		img[2514] = 8'b10011011;
		img[2513] = 8'b10101001;
		img[2512] = 8'b11000001;
		img[2511] = 8'b00101011;
		img[2510] = 8'b00001110;
		img[2509] = 8'b00010010;
		img[2508] = 8'b00100011;
		img[2507] = 8'b00111111;
		img[2506] = 8'b01000111;
		img[2505] = 8'b00100101;
		img[2504] = 8'b00010111;
		img[2503] = 8'b00010000;
		img[2502] = 8'b00010010;
		img[2501] = 8'b00000100;
		img[2500] = 8'b00011000;
		img[2499] = 8'b00000000;
		img[2498] = 8'b00000000;
		img[2497] = 8'b00001110;
		img[2496] = 8'b00000010;
		img[2495] = 8'b00011101;
		img[2494] = 8'b00111101;
		img[2493] = 8'b00100011;
		img[2492] = 8'b00100010;
		img[2491] = 8'b00110010;
		img[2490] = 8'b00001101;
		img[2489] = 8'b00010010;
		img[2488] = 8'b00010101;
		img[2487] = 8'b00001010;
		img[2486] = 8'b00001111;
		img[2485] = 8'b00000110;
		img[2484] = 8'b00001010;
		img[2483] = 8'b00000101;
		img[2482] = 8'b00000101;
		img[2481] = 8'b00001001;
		img[2480] = 8'b00000000;
		img[2479] = 8'b00011100;
		img[2478] = 8'b00000011;
		img[2477] = 8'b00010000;
		img[2476] = 8'b00011111;
		img[2475] = 8'b00110010;
		img[2474] = 8'b00011101;
		img[2473] = 8'b00001111;
		img[2472] = 8'b00000100;
		img[2471] = 8'b00010101;
		img[2470] = 8'b00011001;
		img[2469] = 8'b00010111;
		img[2468] = 8'b00110000;
		img[2467] = 8'b00001111;
		img[2466] = 8'b00001000;
		img[2465] = 8'b00001011;
		img[2464] = 8'b00000000;
		img[2463] = 8'b00100101;
		img[2462] = 8'b00001111;
		img[2461] = 8'b00000000;
		img[2460] = 8'b00101000;
		img[2459] = 8'b00000000;
		img[2458] = 8'b00001010;
		img[2457] = 8'b00011011;
		img[2456] = 8'b00001110;
		img[2455] = 8'b00000100;
		img[2454] = 8'b00001011;
		img[2453] = 8'b00100100;
		img[2452] = 8'b10010100;
		img[2451] = 8'b11000100;
		img[2450] = 8'b10101011;
		img[2449] = 8'b10001100;
		img[2448] = 8'b11001011;
		img[2447] = 8'b10001111;
		img[2446] = 8'b00011001;
		img[2445] = 8'b01000100;
		img[2444] = 8'b01111000;
		img[2443] = 8'b00101100;
		img[2442] = 8'b00101000;
		img[2441] = 8'b00000000;
		img[2440] = 8'b00000010;
		img[2439] = 8'b00001011;
		img[2438] = 8'b00001111;
		img[2437] = 8'b00000101;
		img[2436] = 8'b00000000;
		img[2435] = 8'b00011001;
		img[2434] = 8'b00000000;
		img[2433] = 8'b00000001;
		img[2432] = 8'b00000001;
		img[2431] = 8'b00110011;
		img[2430] = 8'b10000011;
		img[2429] = 8'b00100101;
		img[2428] = 8'b01100101;
		img[2427] = 8'b01000010;
		img[2426] = 8'b00011100;
		img[2425] = 8'b00000000;
		img[2424] = 8'b00100001;
		img[2423] = 8'b00011110;
		img[2422] = 8'b00011010;
		img[2421] = 8'b00101100;
		img[2420] = 8'b00010001;
		img[2419] = 8'b00011011;
		img[2418] = 8'b00001110;
		img[2417] = 8'b00000110;
		img[2416] = 8'b00010010;
		img[2415] = 8'b00000000;
		img[2414] = 8'b00001011;
		img[2413] = 8'b00000000;
		img[2412] = 8'b10000100;
		img[2411] = 8'b01000110;
		img[2410] = 8'b10001011;
		img[2409] = 8'b01101011;
		img[2408] = 8'b01111001;
		img[2407] = 8'b01010101;
		img[2406] = 8'b00010111;
		img[2405] = 8'b00011001;
		img[2404] = 8'b00100110;
		img[2403] = 8'b00010000;
		img[2402] = 8'b00000110;
		img[2401] = 8'b00000000;
		img[2400] = 8'b00001100;
		img[2399] = 8'b00110010;
		img[2398] = 8'b00000000;
		img[2397] = 8'b00010000;
		img[2396] = 8'b00001101;
		img[2395] = 8'b00001110;
		img[2394] = 8'b00010010;
		img[2393] = 8'b00010010;
		img[2392] = 8'b00010011;
		img[2391] = 8'b00011000;
		img[2390] = 8'b00100100;
		img[2389] = 8'b00010100;
		img[2388] = 8'b01011101;
		img[2387] = 8'b01010100;
		img[2386] = 8'b10001011;
		img[2385] = 8'b10100110;
		img[2384] = 8'b10000101;
		img[2383] = 8'b10011010;
		img[2382] = 8'b01011100;
		img[2381] = 8'b01001011;
		img[2380] = 8'b01111111;
		img[2379] = 8'b00001101;
		img[2378] = 8'b00010000;
		img[2377] = 8'b00000000;
		img[2376] = 8'b00000000;
		img[2375] = 8'b00001010;
		img[2374] = 8'b00010110;
		img[2373] = 8'b00010001;
		img[2372] = 8'b00010000;
		img[2371] = 8'b00001100;
		img[2370] = 8'b00001000;
		img[2369] = 8'b00000000;
		img[2368] = 8'b00000000;
		img[2367] = 8'b01100100;
		img[2366] = 8'b10110111;
		img[2365] = 8'b00111001;
		img[2364] = 8'b01111110;
		img[2363] = 8'b01100010;
		img[2362] = 8'b00011101;
		img[2361] = 8'b00001110;
		img[2360] = 8'b00110000;
		img[2359] = 8'b01110011;
		img[2358] = 8'b00011001;
		img[2357] = 8'b00101011;
		img[2356] = 8'b00100110;
		img[2355] = 8'b00011000;
		img[2354] = 8'b00100010;
		img[2353] = 8'b00010101;
		img[2352] = 8'b00000100;
		img[2351] = 8'b00001001;
		img[2350] = 8'b00001010;
		img[2349] = 8'b00010001;
		img[2348] = 8'b00010001;
		img[2347] = 8'b00001001;
		img[2346] = 8'b00101101;
		img[2345] = 8'b01010110;
		img[2344] = 8'b01101001;
		img[2343] = 8'b10000000;
		img[2342] = 8'b00111001;
		img[2341] = 8'b00001001;
		img[2340] = 8'b00000011;
		img[2339] = 8'b00000000;
		img[2338] = 8'b00011110;
		img[2337] = 8'b00000110;
		img[2336] = 8'b00010100;
		img[2335] = 8'b00011100;
		img[2334] = 8'b00010000;
		img[2333] = 8'b00010000;
		img[2332] = 8'b00010001;
		img[2331] = 8'b00010110;
		img[2330] = 8'b00010010;
		img[2329] = 8'b00011011;
		img[2328] = 8'b00011000;
		img[2327] = 8'b00001110;
		img[2326] = 8'b00011111;
		img[2325] = 8'b00000111;
		img[2324] = 8'b00010111;
		img[2323] = 8'b01000101;
		img[2322] = 8'b01101000;
		img[2321] = 8'b10001001;
		img[2320] = 8'b10100110;
		img[2319] = 8'b10111010;
		img[2318] = 8'b10010101;
		img[2317] = 8'b10010000;
		img[2316] = 8'b00111011;
		img[2315] = 8'b00111011;
		img[2314] = 8'b00000001;
		img[2313] = 8'b00010001;
		img[2312] = 8'b00000000;
		img[2311] = 8'b00011010;
		img[2310] = 8'b00001111;
		img[2309] = 8'b00000100;
		img[2308] = 8'b00010000;
		img[2307] = 8'b00001100;
		img[2306] = 8'b00000001;
		img[2305] = 8'b00000101;
		img[2304] = 8'b00001111;
		img[2303] = 8'b01111011;
		img[2302] = 8'b10001011;
		img[2301] = 8'b01000101;
		img[2300] = 8'b01011101;
		img[2299] = 8'b00100011;
		img[2298] = 8'b00101111;
		img[2297] = 8'b00101011;
		img[2296] = 8'b01011011;
		img[2295] = 8'b01000100;
		img[2294] = 8'b00011010;
		img[2293] = 8'b00101100;
		img[2292] = 8'b00101110;
		img[2291] = 8'b00100000;
		img[2290] = 8'b00100010;
		img[2289] = 8'b00100001;
		img[2288] = 8'b00011101;
		img[2287] = 8'b00100101;
		img[2286] = 8'b00010100;
		img[2285] = 8'b00001101;
		img[2284] = 8'b00010000;
		img[2283] = 8'b00000000;
		img[2282] = 8'b00010010;
		img[2281] = 8'b00000001;
		img[2280] = 8'b01000000;
		img[2279] = 8'b00110110;
		img[2278] = 8'b01111100;
		img[2277] = 8'b00001101;
		img[2276] = 8'b00100110;
		img[2275] = 8'b00000001;
		img[2274] = 8'b00011110;
		img[2273] = 8'b00001110;
		img[2272] = 8'b00010001;
		img[2271] = 8'b00011000;
		img[2270] = 8'b00010101;
		img[2269] = 8'b00001011;
		img[2268] = 8'b00010010;
		img[2267] = 8'b00001100;
		img[2266] = 8'b00010111;
		img[2265] = 8'b00011010;
		img[2264] = 8'b00100010;
		img[2263] = 8'b00001100;
		img[2262] = 8'b00001110;
		img[2261] = 8'b00010000;
		img[2260] = 8'b00000011;
		img[2259] = 8'b10011101;
		img[2258] = 8'b11000010;
		img[2257] = 8'b11001010;
		img[2256] = 8'b10010111;
		img[2255] = 8'b10000110;
		img[2254] = 8'b10100100;
		img[2253] = 8'b01100011;
		img[2252] = 8'b01110111;
		img[2251] = 8'b00100110;
		img[2250] = 8'b00000000;
		img[2249] = 8'b00000101;
		img[2248] = 8'b00000100;
		img[2247] = 8'b00000100;
		img[2246] = 8'b00001110;
		img[2245] = 8'b00010100;
		img[2244] = 8'b00010011;
		img[2243] = 8'b00010010;
		img[2242] = 8'b00001101;
		img[2241] = 8'b00010110;
		img[2240] = 8'b00000000;
		img[2239] = 8'b01010110;
		img[2238] = 8'b01100000;
		img[2237] = 8'b00111000;
		img[2236] = 8'b01111010;
		img[2235] = 8'b10001111;
		img[2234] = 8'b00011101;
		img[2233] = 8'b01101011;
		img[2232] = 8'b01011101;
		img[2231] = 8'b00111100;
		img[2230] = 8'b00101101;
		img[2229] = 8'b00100000;
		img[2228] = 8'b00010100;
		img[2227] = 8'b00011010;
		img[2226] = 8'b00011011;
		img[2225] = 8'b00011000;
		img[2224] = 8'b00011000;
		img[2223] = 8'b00110011;
		img[2222] = 8'b00011101;
		img[2221] = 8'b00011100;
		img[2220] = 8'b00001100;
		img[2219] = 8'b00001100;
		img[2218] = 8'b00011011;
		img[2217] = 8'b00001110;
		img[2216] = 8'b00001101;
		img[2215] = 8'b00001100;
		img[2214] = 8'b00111000;
		img[2213] = 8'b00101110;
		img[2212] = 8'b00011001;
		img[2211] = 8'b00010100;
		img[2210] = 8'b00101011;
		img[2209] = 8'b00000100;
		img[2208] = 8'b00001100;
		img[2207] = 8'b00000101;
		img[2206] = 8'b00010110;
		img[2205] = 8'b00011010;
		img[2204] = 8'b00010011;
		img[2203] = 8'b00100011;
		img[2202] = 8'b00101001;
		img[2201] = 8'b00011111;
		img[2200] = 8'b00010101;
		img[2199] = 8'b00010101;
		img[2198] = 8'b00010011;
		img[2197] = 8'b00001011;
		img[2196] = 8'b00010000;
		img[2195] = 8'b00001101;
		img[2194] = 8'b00110111;
		img[2193] = 8'b11001011;
		img[2192] = 8'b11100001;
		img[2191] = 8'b10111100;
		img[2190] = 8'b10110011;
		img[2189] = 8'b10011100;
		img[2188] = 8'b10001111;
		img[2187] = 8'b00101011;
		img[2186] = 8'b00100010;
		img[2185] = 8'b00000000;
		img[2184] = 8'b00001100;
		img[2183] = 8'b00000000;
		img[2182] = 8'b00010111;
		img[2181] = 8'b00001111;
		img[2180] = 8'b00001100;
		img[2179] = 8'b00010001;
		img[2178] = 8'b00001111;
		img[2177] = 8'b00001100;
		img[2176] = 8'b00000000;
		img[2175] = 8'b00111011;
		img[2174] = 8'b01000011;
		img[2173] = 8'b01101011;
		img[2172] = 8'b10010101;
		img[2171] = 8'b00110111;
		img[2170] = 8'b01111101;
		img[2169] = 8'b01101000;
		img[2168] = 8'b01001011;
		img[2167] = 8'b00110010;
		img[2166] = 8'b00111000;
		img[2165] = 8'b00100011;
		img[2164] = 8'b00111011;
		img[2163] = 8'b00100100;
		img[2162] = 8'b00101100;
		img[2161] = 8'b00011101;
		img[2160] = 8'b00100000;
		img[2159] = 8'b00010111;
		img[2158] = 8'b00101010;
		img[2157] = 8'b00110011;
		img[2156] = 8'b00110111;
		img[2155] = 8'b00001101;
		img[2154] = 8'b00001000;
		img[2153] = 8'b00000100;
		img[2152] = 8'b00011001;
		img[2151] = 8'b00100111;
		img[2150] = 8'b01100001;
		img[2149] = 8'b01000001;
		img[2148] = 8'b00100001;
		img[2147] = 8'b00000101;
		img[2146] = 8'b00010001;
		img[2145] = 8'b00011100;
		img[2144] = 8'b00100111;
		img[2143] = 8'b00001001;
		img[2142] = 8'b00100011;
		img[2141] = 8'b00100101;
		img[2140] = 8'b00010001;
		img[2139] = 8'b01100010;
		img[2138] = 8'b00110101;
		img[2137] = 8'b01000110;
		img[2136] = 8'b01010100;
		img[2135] = 8'b00011101;
		img[2134] = 8'b00101001;
		img[2133] = 8'b00100011;
		img[2132] = 8'b00011100;
		img[2131] = 8'b00011010;
		img[2130] = 8'b00100111;
		img[2129] = 8'b01010100;
		img[2128] = 8'b01000111;
		img[2127] = 8'b00101101;
		img[2126] = 8'b00111010;
		img[2125] = 8'b01101011;
		img[2124] = 8'b01010010;
		img[2123] = 8'b00100100;
		img[2122] = 8'b00011001;
		img[2121] = 8'b00001000;
		img[2120] = 8'b00010001;
		img[2119] = 8'b00001101;
		img[2118] = 8'b00000111;
		img[2117] = 8'b00000010;
		img[2116] = 8'b00000101;
		img[2115] = 8'b00001010;
		img[2114] = 8'b00001100;
		img[2113] = 8'b00001011;
		img[2112] = 8'b00000000;
		img[2111] = 8'b01100010;
		img[2110] = 8'b10000010;
		img[2109] = 8'b10001000;
		img[2108] = 8'b01011010;
		img[2107] = 8'b10110000;
		img[2106] = 8'b01100100;
		img[2105] = 8'b01111100;
		img[2104] = 8'b01010000;
		img[2103] = 8'b01110010;
		img[2102] = 8'b01101110;
		img[2101] = 8'b00110111;
		img[2100] = 8'b01010001;
		img[2099] = 8'b00101001;
		img[2098] = 8'b00100101;
		img[2097] = 8'b01000000;
		img[2096] = 8'b00111000;
		img[2095] = 8'b00001101;
		img[2094] = 8'b00111001;
		img[2093] = 8'b10000001;
		img[2092] = 8'b00110001;
		img[2091] = 8'b00100000;
		img[2090] = 8'b00011010;
		img[2089] = 8'b00101010;
		img[2088] = 8'b00010111;
		img[2087] = 8'b01000100;
		img[2086] = 8'b10011111;
		img[2085] = 8'b11001101;
		img[2084] = 8'b10011111;
		img[2083] = 8'b01000100;
		img[2082] = 8'b00011000;
		img[2081] = 8'b00001111;
		img[2080] = 8'b00011101;
		img[2079] = 8'b00010101;
		img[2078] = 8'b00101110;
		img[2077] = 8'b00100101;
		img[2076] = 8'b01001111;
		img[2075] = 8'b01010100;
		img[2074] = 8'b01101000;
		img[2073] = 8'b10100001;
		img[2072] = 8'b01011110;
		img[2071] = 8'b01000010;
		img[2070] = 8'b00100110;
		img[2069] = 8'b00101010;
		img[2068] = 8'b00100001;
		img[2067] = 8'b00010001;
		img[2066] = 8'b01001010;
		img[2065] = 8'b01010100;
		img[2064] = 8'b01000111;
		img[2063] = 8'b00111011;
		img[2062] = 8'b01000111;
		img[2061] = 8'b01111001;
		img[2060] = 8'b01111110;
		img[2059] = 8'b01011000;
		img[2058] = 8'b00000111;
		img[2057] = 8'b00010111;
		img[2056] = 8'b00001010;
		img[2055] = 8'b00010000;
		img[2054] = 8'b00010011;
		img[2053] = 8'b00001011;
		img[2052] = 8'b00001010;
		img[2051] = 8'b00001010;
		img[2050] = 8'b00001101;
		img[2049] = 8'b00000000;
		img[2048] = 8'b00000000;
		img[2047] = 8'b10011001;
		img[2046] = 8'b10000101;
		img[2045] = 8'b01011010;
		img[2044] = 8'b01101001;
		img[2043] = 8'b10111111;
		img[2042] = 8'b01110010;
		img[2041] = 8'b01011011;
		img[2040] = 8'b01111000;
		img[2039] = 8'b01011000;
		img[2038] = 8'b01110101;
		img[2037] = 8'b10000001;
		img[2036] = 8'b01101101;
		img[2035] = 8'b01000110;
		img[2034] = 8'b01100011;
		img[2033] = 8'b00101100;
		img[2032] = 8'b01010010;
		img[2031] = 8'b00101001;
		img[2030] = 8'b01011110;
		img[2029] = 8'b01110110;
		img[2028] = 8'b00110110;
		img[2027] = 8'b00100101;
		img[2026] = 8'b00101111;
		img[2025] = 8'b00111110;
		img[2024] = 8'b00100001;
		img[2023] = 8'b00011010;
		img[2022] = 8'b01010000;
		img[2021] = 8'b10001110;
		img[2020] = 8'b10110001;
		img[2019] = 8'b11100110;
		img[2018] = 8'b10011001;
		img[2017] = 8'b01001010;
		img[2016] = 8'b01001000;
		img[2015] = 8'b01100011;
		img[2014] = 8'b01100010;
		img[2013] = 8'b01111101;
		img[2012] = 8'b01110001;
		img[2011] = 8'b10010101;
		img[2010] = 8'b10101100;
		img[2009] = 8'b11001000;
		img[2008] = 8'b10011111;
		img[2007] = 8'b10010110;
		img[2006] = 8'b01101001;
		img[2005] = 8'b01000101;
		img[2004] = 8'b01001111;
		img[2003] = 8'b01101110;
		img[2002] = 8'b01110111;
		img[2001] = 8'b10011101;
		img[2000] = 8'b10001000;
		img[1999] = 8'b01111111;
		img[1998] = 8'b10000001;
		img[1997] = 8'b10001000;
		img[1996] = 8'b01111101;
		img[1995] = 8'b01101110;
		img[1994] = 8'b01001100;
		img[1993] = 8'b00011111;
		img[1992] = 8'b00101100;
		img[1991] = 8'b00001011;
		img[1990] = 8'b00000000;
		img[1989] = 8'b00000000;
		img[1988] = 8'b00100011;
		img[1987] = 8'b00000111;
		img[1986] = 8'b00000010;
		img[1985] = 8'b00001011;
		img[1984] = 8'b00000110;
		img[1983] = 8'b01001010;
		img[1982] = 8'b00110001;
		img[1981] = 8'b01101100;
		img[1980] = 8'b01010011;
		img[1979] = 8'b01101100;
		img[1978] = 8'b01011111;
		img[1977] = 8'b01011001;
		img[1976] = 8'b01010011;
		img[1975] = 8'b01110110;
		img[1974] = 8'b01011010;
		img[1973] = 8'b01100000;
		img[1972] = 8'b10000110;
		img[1971] = 8'b00001110;
		img[1970] = 8'b00111000;
		img[1969] = 8'b01000000;
		img[1968] = 8'b01100000;
		img[1967] = 8'b01100011;
		img[1966] = 8'b01110010;
		img[1965] = 8'b01010001;
		img[1964] = 8'b01110110;
		img[1963] = 8'b00011001;
		img[1962] = 8'b00001101;
		img[1961] = 8'b00010101;
		img[1960] = 8'b00111001;
		img[1959] = 8'b01000000;
		img[1958] = 8'b10001110;
		img[1957] = 8'b10111101;
		img[1956] = 8'b10111110;
		img[1955] = 8'b11010000;
		img[1954] = 8'b11000110;
		img[1953] = 8'b01110000;
		img[1952] = 8'b10011000;
		img[1951] = 8'b10001101;
		img[1950] = 8'b10100100;
		img[1949] = 8'b01111010;
		img[1948] = 8'b10001000;
		img[1947] = 8'b01111001;
		img[1946] = 8'b10101001;
		img[1945] = 8'b10010110;
		img[1944] = 8'b01111000;
		img[1943] = 8'b10000011;
		img[1942] = 8'b01100011;
		img[1941] = 8'b10001011;
		img[1940] = 8'b01110110;
		img[1939] = 8'b01101100;
		img[1938] = 8'b10001100;
		img[1937] = 8'b10001101;
		img[1936] = 8'b10001001;
		img[1935] = 8'b10001100;
		img[1934] = 8'b10001010;
		img[1933] = 8'b01110100;
		img[1932] = 8'b01110000;
		img[1931] = 8'b01011100;
		img[1930] = 8'b01011101;
		img[1929] = 8'b00110111;
		img[1928] = 8'b01010000;
		img[1927] = 8'b00101101;
		img[1926] = 8'b00010010;
		img[1925] = 8'b00000000;
		img[1924] = 8'b00010111;
		img[1923] = 8'b00001100;
		img[1922] = 8'b00000000;
		img[1921] = 8'b00000000;
		img[1920] = 8'b00000110;
		img[1919] = 8'b01110110;
		img[1918] = 8'b10000100;
		img[1917] = 8'b10000011;
		img[1916] = 8'b10010010;
		img[1915] = 8'b01101011;
		img[1914] = 8'b01110010;
		img[1913] = 8'b01111111;
		img[1912] = 8'b01100110;
		img[1911] = 8'b10001010;
		img[1910] = 8'b01101110;
		img[1909] = 8'b10001001;
		img[1908] = 8'b10001110;
		img[1907] = 8'b01101010;
		img[1906] = 8'b10101000;
		img[1905] = 8'b10111100;
		img[1904] = 8'b10101010;
		img[1903] = 8'b10111110;
		img[1902] = 8'b10101000;
		img[1901] = 8'b10111111;
		img[1900] = 8'b11000101;
		img[1899] = 8'b01110001;
		img[1898] = 8'b10010001;
		img[1897] = 8'b00110110;
		img[1896] = 8'b01111010;
		img[1895] = 8'b11000010;
		img[1894] = 8'b10101110;
		img[1893] = 8'b10011110;
		img[1892] = 8'b10010101;
		img[1891] = 8'b10100000;
		img[1890] = 8'b10010011;
		img[1889] = 8'b10110001;
		img[1888] = 8'b10101011;
		img[1887] = 8'b10011111;
		img[1886] = 8'b10101000;
		img[1885] = 8'b01111101;
		img[1884] = 8'b10000111;
		img[1883] = 8'b11010101;
		img[1882] = 8'b10011001;
		img[1881] = 8'b10101101;
		img[1880] = 8'b10011001;
		img[1879] = 8'b10000001;
		img[1878] = 8'b01111110;
		img[1877] = 8'b10000001;
		img[1876] = 8'b10010010;
		img[1875] = 8'b10110010;
		img[1874] = 8'b10000111;
		img[1873] = 8'b01001000;
		img[1872] = 8'b01000000;
		img[1871] = 8'b00101001;
		img[1870] = 8'b00111101;
		img[1869] = 8'b01110110;
		img[1868] = 8'b00110010;
		img[1867] = 8'b00111001;
		img[1866] = 8'b00111011;
		img[1865] = 8'b00100011;
		img[1864] = 8'b00100001;
		img[1863] = 8'b00000000;
		img[1862] = 8'b00001010;
		img[1861] = 8'b00010000;
		img[1860] = 8'b00010001;
		img[1859] = 8'b00000110;
		img[1858] = 8'b00001000;
		img[1857] = 8'b00000000;
		img[1856] = 8'b00000100;
		img[1855] = 8'b01110011;
		img[1854] = 8'b01100101;
		img[1853] = 8'b01101001;
		img[1852] = 8'b10010010;
		img[1851] = 8'b01101101;
		img[1850] = 8'b01111101;
		img[1849] = 8'b01111011;
		img[1848] = 8'b10010101;
		img[1847] = 8'b10111111;
		img[1846] = 8'b10100100;
		img[1845] = 8'b10011110;
		img[1844] = 8'b10110000;
		img[1843] = 8'b10011010;
		img[1842] = 8'b10101110;
		img[1841] = 8'b11010110;
		img[1840] = 8'b11011110;
		img[1839] = 8'b11110001;
		img[1838] = 8'b11110110;
		img[1837] = 8'b11100100;
		img[1836] = 8'b11010001;
		img[1835] = 8'b11010000;
		img[1834] = 8'b11011000;
		img[1833] = 8'b10101110;
		img[1832] = 8'b11010011;
		img[1831] = 8'b11010010;
		img[1830] = 8'b11100010;
		img[1829] = 8'b11101100;
		img[1828] = 8'b11101011;
		img[1827] = 8'b11100001;
		img[1826] = 8'b11100011;
		img[1825] = 8'b11100010;
		img[1824] = 8'b11010000;
		img[1823] = 8'b11010110;
		img[1822] = 8'b10111111;
		img[1821] = 8'b10110111;
		img[1820] = 8'b10011110;
		img[1819] = 8'b10011110;
		img[1818] = 8'b10110001;
		img[1817] = 8'b10010010;
		img[1816] = 8'b01111100;
		img[1815] = 8'b01011001;
		img[1814] = 8'b01001110;
		img[1813] = 8'b01010110;
		img[1812] = 8'b01000100;
		img[1811] = 8'b01011101;
		img[1810] = 8'b01010101;
		img[1809] = 8'b00011110;
		img[1808] = 8'b00010101;
		img[1807] = 8'b00000110;
		img[1806] = 8'b00010000;
		img[1805] = 8'b01011010;
		img[1804] = 8'b00101101;
		img[1803] = 8'b00100011;
		img[1802] = 8'b00101110;
		img[1801] = 8'b00011011;
		img[1800] = 8'b00011100;
		img[1799] = 8'b00000001;
		img[1798] = 8'b00000100;
		img[1797] = 8'b00000000;
		img[1796] = 8'b00010111;
		img[1795] = 8'b00001010;
		img[1794] = 8'b00011110;
		img[1793] = 8'b00001110;
		img[1792] = 8'b00000000;
		img[1791] = 8'b01000011;
		img[1790] = 8'b01001100;
		img[1789] = 8'b00111111;
		img[1788] = 8'b01001111;
		img[1787] = 8'b01010001;
		img[1786] = 8'b01100001;
		img[1785] = 8'b01100110;
		img[1784] = 8'b01100111;
		img[1783] = 8'b10001101;
		img[1782] = 8'b10100100;
		img[1781] = 8'b11000110;
		img[1780] = 8'b10100010;
		img[1779] = 8'b11001011;
		img[1778] = 8'b10100100;
		img[1777] = 8'b11010011;
		img[1776] = 8'b11100010;
		img[1775] = 8'b11011110;
		img[1774] = 8'b11011001;
		img[1773] = 8'b11000001;
		img[1772] = 8'b11010110;
		img[1771] = 8'b10111111;
		img[1770] = 8'b10100010;
		img[1769] = 8'b10111000;
		img[1768] = 8'b10011101;
		img[1767] = 8'b10100011;
		img[1766] = 8'b10101110;
		img[1765] = 8'b10111011;
		img[1764] = 8'b11010001;
		img[1763] = 8'b11000101;
		img[1762] = 8'b10111010;
		img[1761] = 8'b11000000;
		img[1760] = 8'b10100010;
		img[1759] = 8'b10011100;
		img[1758] = 8'b10110001;
		img[1757] = 8'b10001111;
		img[1756] = 8'b01110111;
		img[1755] = 8'b01110001;
		img[1754] = 8'b10000001;
		img[1753] = 8'b10000011;
		img[1752] = 8'b01110111;
		img[1751] = 8'b01010000;
		img[1750] = 8'b01001000;
		img[1749] = 8'b01001101;
		img[1748] = 8'b00110010;
		img[1747] = 8'b01011100;
		img[1746] = 8'b01010101;
		img[1745] = 8'b00010110;
		img[1744] = 8'b00000111;
		img[1743] = 8'b00000000;
		img[1742] = 8'b00000000;
		img[1741] = 8'b01011010;
		img[1740] = 8'b00100101;
		img[1739] = 8'b00011001;
		img[1738] = 8'b00111111;
		img[1737] = 8'b00001111;
		img[1736] = 8'b00010100;
		img[1735] = 8'b00001011;
		img[1734] = 8'b00000111;
		img[1733] = 8'b00000111;
		img[1732] = 8'b00001110;
		img[1731] = 8'b00000110;
		img[1730] = 8'b00000000;
		img[1729] = 8'b00011100;
		img[1728] = 8'b00001110;
		img[1727] = 8'b00110000;
		img[1726] = 8'b00110010;
		img[1725] = 8'b01001000;
		img[1724] = 8'b01001011;
		img[1723] = 8'b00111010;
		img[1722] = 8'b01010001;
		img[1721] = 8'b01011101;
		img[1720] = 8'b01101011;
		img[1719] = 8'b01111101;
		img[1718] = 8'b10010100;
		img[1717] = 8'b10101100;
		img[1716] = 8'b10111011;
		img[1715] = 8'b11000000;
		img[1714] = 8'b11000100;
		img[1713] = 8'b11001101;
		img[1712] = 8'b11010110;
		img[1711] = 8'b11001111;
		img[1710] = 8'b11000011;
		img[1709] = 8'b10101011;
		img[1708] = 8'b11000011;
		img[1707] = 8'b10011011;
		img[1706] = 8'b10001101;
		img[1705] = 8'b10100111;
		img[1704] = 8'b01110011;
		img[1703] = 8'b01110111;
		img[1702] = 8'b01111101;
		img[1701] = 8'b10000101;
		img[1700] = 8'b11000011;
		img[1699] = 8'b11000100;
		img[1698] = 8'b10110001;
		img[1697] = 8'b10110000;
		img[1696] = 8'b01111010;
		img[1695] = 8'b10001100;
		img[1694] = 8'b10101001;
		img[1693] = 8'b01100010;
		img[1692] = 8'b01011011;
		img[1691] = 8'b01111011;
		img[1690] = 8'b01101100;
		img[1689] = 8'b01111111;
		img[1688] = 8'b01101101;
		img[1687] = 8'b01001111;
		img[1686] = 8'b01000110;
		img[1685] = 8'b01001101;
		img[1684] = 8'b00100011;
		img[1683] = 8'b01010101;
		img[1682] = 8'b01100000;
		img[1681] = 8'b00010100;
		img[1680] = 8'b00000111;
		img[1679] = 8'b00000000;
		img[1678] = 8'b00001000;
		img[1677] = 8'b01001000;
		img[1676] = 8'b00101111;
		img[1675] = 8'b00010110;
		img[1674] = 8'b00111001;
		img[1673] = 8'b00001001;
		img[1672] = 8'b00011101;
		img[1671] = 8'b00001010;
		img[1670] = 8'b00011000;
		img[1669] = 8'b00011011;
		img[1668] = 8'b00001110;
		img[1667] = 8'b00000001;
		img[1666] = 8'b00001110;
		img[1665] = 8'b00000000;
		img[1664] = 8'b00011110;
		img[1663] = 8'b00100111;
		img[1662] = 8'b00110101;
		img[1661] = 8'b00111100;
		img[1660] = 8'b01000010;
		img[1659] = 8'b01000110;
		img[1658] = 8'b01000101;
		img[1657] = 8'b01010011;
		img[1656] = 8'b01100010;
		img[1655] = 8'b01110111;
		img[1654] = 8'b10000000;
		img[1653] = 8'b10100000;
		img[1652] = 8'b10110010;
		img[1651] = 8'b10011100;
		img[1650] = 8'b11010000;
		img[1649] = 8'b11001010;
		img[1648] = 8'b11010001;
		img[1647] = 8'b11010011;
		img[1646] = 8'b10111101;
		img[1645] = 8'b10110101;
		img[1644] = 8'b10111010;
		img[1643] = 8'b10011010;
		img[1642] = 8'b10010010;
		img[1641] = 8'b10011111;
		img[1640] = 8'b01100100;
		img[1639] = 8'b01011011;
		img[1638] = 8'b01001011;
		img[1637] = 8'b01010011;
		img[1636] = 8'b10100110;
		img[1635] = 8'b11001101;
		img[1634] = 8'b10100110;
		img[1633] = 8'b10101011;
		img[1632] = 8'b01011100;
		img[1631] = 8'b01111100;
		img[1630] = 8'b10101111;
		img[1629] = 8'b10000111;
		img[1628] = 8'b00111111;
		img[1627] = 8'b01110000;
		img[1626] = 8'b01110001;
		img[1625] = 8'b10010010;
		img[1624] = 8'b01101000;
		img[1623] = 8'b01001011;
		img[1622] = 8'b01000110;
		img[1621] = 8'b01010000;
		img[1620] = 8'b00100000;
		img[1619] = 8'b01011000;
		img[1618] = 8'b01100111;
		img[1617] = 8'b00010001;
		img[1616] = 8'b00001100;
		img[1615] = 8'b00000011;
		img[1614] = 8'b00000001;
		img[1613] = 8'b01000001;
		img[1612] = 8'b00110011;
		img[1611] = 8'b00010110;
		img[1610] = 8'b00110100;
		img[1609] = 8'b00010000;
		img[1608] = 8'b00100000;
		img[1607] = 8'b00010001;
		img[1606] = 8'b00010111;
		img[1605] = 8'b00011001;
		img[1604] = 8'b00100011;
		img[1603] = 8'b00010111;
		img[1602] = 8'b00001111;
		img[1601] = 8'b00001100;
		img[1600] = 8'b00000110;
		img[1599] = 8'b00101001;
		img[1598] = 8'b00100111;
		img[1597] = 8'b00101001;
		img[1596] = 8'b00111001;
		img[1595] = 8'b00111100;
		img[1594] = 8'b00111011;
		img[1593] = 8'b01000100;
		img[1592] = 8'b01011011;
		img[1591] = 8'b01100111;
		img[1590] = 8'b01111010;
		img[1589] = 8'b10000110;
		img[1588] = 8'b10111010;
		img[1587] = 8'b11000010;
		img[1586] = 8'b10111111;
		img[1585] = 8'b11000111;
		img[1584] = 8'b11010010;
		img[1583] = 8'b11011000;
		img[1582] = 8'b11001001;
		img[1581] = 8'b11001101;
		img[1580] = 8'b10110100;
		img[1579] = 8'b10100000;
		img[1578] = 8'b10001100;
		img[1577] = 8'b10001101;
		img[1576] = 8'b01101010;
		img[1575] = 8'b01010110;
		img[1574] = 8'b00110100;
		img[1573] = 8'b00111001;
		img[1572] = 8'b10001011;
		img[1571] = 8'b11010000;
		img[1570] = 8'b10101100;
		img[1569] = 8'b10101101;
		img[1568] = 8'b01010000;
		img[1567] = 8'b01111001;
		img[1566] = 8'b10101111;
		img[1565] = 8'b01111000;
		img[1564] = 8'b01010100;
		img[1563] = 8'b01110001;
		img[1562] = 8'b01100100;
		img[1561] = 8'b10010100;
		img[1560] = 8'b01100100;
		img[1559] = 8'b01001001;
		img[1558] = 8'b01000011;
		img[1557] = 8'b01010000;
		img[1556] = 8'b00011011;
		img[1555] = 8'b01010011;
		img[1554] = 8'b01110000;
		img[1553] = 8'b00010000;
		img[1552] = 8'b00001011;
		img[1551] = 8'b00000000;
		img[1550] = 8'b00000010;
		img[1549] = 8'b01000100;
		img[1548] = 8'b01000110;
		img[1547] = 8'b00011001;
		img[1546] = 8'b00101101;
		img[1545] = 8'b00100111;
		img[1544] = 8'b00100001;
		img[1543] = 8'b00010010;
		img[1542] = 8'b00011111;
		img[1541] = 8'b00011101;
		img[1540] = 8'b00000101;
		img[1539] = 8'b00100000;
		img[1538] = 8'b00001110;
		img[1537] = 8'b00000000;
		img[1536] = 8'b00000000;
		img[1535] = 8'b00010011;
		img[1534] = 8'b00011101;
		img[1533] = 8'b00100111;
		img[1532] = 8'b00110111;
		img[1531] = 8'b00101011;
		img[1530] = 8'b00110000;
		img[1529] = 8'b00111100;
		img[1528] = 8'b01001000;
		img[1527] = 8'b01010101;
		img[1526] = 8'b01101100;
		img[1525] = 8'b01110011;
		img[1524] = 8'b10100100;
		img[1523] = 8'b10111010;
		img[1522] = 8'b10111010;
		img[1521] = 8'b11001010;
		img[1520] = 8'b11001101;
		img[1519] = 8'b11010110;
		img[1518] = 8'b11001110;
		img[1517] = 8'b11011000;
		img[1516] = 8'b10100111;
		img[1515] = 8'b10110010;
		img[1514] = 8'b10001111;
		img[1513] = 8'b10000011;
		img[1512] = 8'b01110010;
		img[1511] = 8'b01011000;
		img[1510] = 8'b00101101;
		img[1509] = 8'b00100101;
		img[1508] = 8'b01101111;
		img[1507] = 8'b11001000;
		img[1506] = 8'b10110111;
		img[1505] = 8'b10110011;
		img[1504] = 8'b01010000;
		img[1503] = 8'b01110100;
		img[1502] = 8'b10100001;
		img[1501] = 8'b01111100;
		img[1500] = 8'b01100010;
		img[1499] = 8'b01110010;
		img[1498] = 8'b01100110;
		img[1497] = 8'b10001100;
		img[1496] = 8'b01100101;
		img[1495] = 8'b01000011;
		img[1494] = 8'b00111101;
		img[1493] = 8'b01010011;
		img[1492] = 8'b00011100;
		img[1491] = 8'b01011011;
		img[1490] = 8'b10000001;
		img[1489] = 8'b00010101;
		img[1488] = 8'b00010001;
		img[1487] = 8'b00001101;
		img[1486] = 8'b00001000;
		img[1485] = 8'b00111011;
		img[1484] = 8'b01011011;
		img[1483] = 8'b00011001;
		img[1482] = 8'b00110000;
		img[1481] = 8'b00001110;
		img[1480] = 8'b00110111;
		img[1479] = 8'b00100111;
		img[1478] = 8'b00000101;
		img[1477] = 8'b00110000;
		img[1476] = 8'b00001011;
		img[1475] = 8'b00100000;
		img[1474] = 8'b00001100;
		img[1473] = 8'b00100000;
		img[1472] = 8'b00011010;
		img[1471] = 8'b00001111;
		img[1470] = 8'b00010101;
		img[1469] = 8'b00100101;
		img[1468] = 8'b00100011;
		img[1467] = 8'b00011011;
		img[1466] = 8'b00110101;
		img[1465] = 8'b00100010;
		img[1464] = 8'b00110100;
		img[1463] = 8'b01001010;
		img[1462] = 8'b01011101;
		img[1461] = 8'b01110010;
		img[1460] = 8'b10000110;
		img[1459] = 8'b10100101;
		img[1458] = 8'b10111001;
		img[1457] = 8'b11000100;
		img[1456] = 8'b11001110;
		img[1455] = 8'b11010001;
		img[1454] = 8'b11010111;
		img[1453] = 8'b11001001;
		img[1452] = 8'b10101111;
		img[1451] = 8'b11000110;
		img[1450] = 8'b10001010;
		img[1449] = 8'b10000011;
		img[1448] = 8'b10001001;
		img[1447] = 8'b01011001;
		img[1446] = 8'b00101010;
		img[1445] = 8'b00011010;
		img[1444] = 8'b01010101;
		img[1443] = 8'b11010100;
		img[1442] = 8'b10111100;
		img[1441] = 8'b10111101;
		img[1440] = 8'b01011101;
		img[1439] = 8'b01110000;
		img[1438] = 8'b10011001;
		img[1437] = 8'b01111000;
		img[1436] = 8'b01111001;
		img[1435] = 8'b01110110;
		img[1434] = 8'b01101001;
		img[1433] = 8'b10000010;
		img[1432] = 8'b01100110;
		img[1431] = 8'b01000000;
		img[1430] = 8'b00111010;
		img[1429] = 8'b01011011;
		img[1428] = 8'b00011111;
		img[1427] = 8'b01100101;
		img[1426] = 8'b10001110;
		img[1425] = 8'b00011101;
		img[1424] = 8'b00000110;
		img[1423] = 8'b00001100;
		img[1422] = 8'b00000100;
		img[1421] = 8'b00101101;
		img[1420] = 8'b01110100;
		img[1419] = 8'b00010011;
		img[1418] = 8'b00011011;
		img[1417] = 8'b00011001;
		img[1416] = 8'b00100010;
		img[1415] = 8'b00010000;
		img[1414] = 8'b00100010;
		img[1413] = 8'b01010000;
		img[1412] = 8'b00011010;
		img[1411] = 8'b00101100;
		img[1410] = 8'b00101100;
		img[1409] = 8'b00000010;
		img[1408] = 8'b00101000;
		img[1407] = 8'b00011100;
		img[1406] = 8'b00010111;
		img[1405] = 8'b00001100;
		img[1404] = 8'b00011101;
		img[1403] = 8'b00011000;
		img[1402] = 8'b00011100;
		img[1401] = 8'b00101100;
		img[1400] = 8'b00110100;
		img[1399] = 8'b01000110;
		img[1398] = 8'b01000110;
		img[1397] = 8'b01111011;
		img[1396] = 8'b01111011;
		img[1395] = 8'b10011001;
		img[1394] = 8'b10110100;
		img[1393] = 8'b10111011;
		img[1392] = 8'b11001011;
		img[1391] = 8'b11011001;
		img[1390] = 8'b11001010;
		img[1389] = 8'b11001000;
		img[1388] = 8'b11000010;
		img[1387] = 8'b11011000;
		img[1386] = 8'b10010011;
		img[1385] = 8'b10000110;
		img[1384] = 8'b10011000;
		img[1383] = 8'b01010010;
		img[1382] = 8'b00011010;
		img[1381] = 8'b00010000;
		img[1380] = 8'b01000010;
		img[1379] = 8'b11011110;
		img[1378] = 8'b10111100;
		img[1377] = 8'b11001100;
		img[1376] = 8'b01101110;
		img[1375] = 8'b01011100;
		img[1374] = 8'b10000011;
		img[1373] = 8'b10000101;
		img[1372] = 8'b10001010;
		img[1371] = 8'b01111111;
		img[1370] = 8'b01101000;
		img[1369] = 8'b01110011;
		img[1368] = 8'b01101011;
		img[1367] = 8'b00110101;
		img[1366] = 8'b00111001;
		img[1365] = 8'b01011001;
		img[1364] = 8'b00010110;
		img[1363] = 8'b01110101;
		img[1362] = 8'b10100100;
		img[1361] = 8'b00111001;
		img[1360] = 8'b00000111;
		img[1359] = 8'b00000000;
		img[1358] = 8'b00010110;
		img[1357] = 8'b00100111;
		img[1356] = 8'b01111110;
		img[1355] = 8'b00011100;
		img[1354] = 8'b00110010;
		img[1353] = 8'b00011001;
		img[1352] = 8'b00011101;
		img[1351] = 8'b00001010;
		img[1350] = 8'b00011111;
		img[1349] = 8'b00111000;
		img[1348] = 8'b00100001;
		img[1347] = 8'b00011000;
		img[1346] = 8'b00001000;
		img[1345] = 8'b00011110;
		img[1344] = 8'b00100000;
		img[1343] = 8'b00001111;
		img[1342] = 8'b00001001;
		img[1341] = 8'b00001100;
		img[1340] = 8'b00000111;
		img[1339] = 8'b00011101;
		img[1338] = 8'b00011011;
		img[1337] = 8'b00100100;
		img[1336] = 8'b00110100;
		img[1335] = 8'b01000011;
		img[1334] = 8'b01011111;
		img[1333] = 8'b01110010;
		img[1332] = 8'b01110011;
		img[1331] = 8'b10001000;
		img[1330] = 8'b10110011;
		img[1329] = 8'b11000100;
		img[1328] = 8'b11001101;
		img[1327] = 8'b11011011;
		img[1326] = 8'b11000110;
		img[1325] = 8'b11001011;
		img[1324] = 8'b11101000;
		img[1323] = 8'b11001010;
		img[1322] = 8'b10110010;
		img[1321] = 8'b10000110;
		img[1320] = 8'b10110010;
		img[1319] = 8'b01010100;
		img[1318] = 8'b00010011;
		img[1317] = 8'b00000110;
		img[1316] = 8'b00100111;
		img[1315] = 8'b11100101;
		img[1314] = 8'b11010000;
		img[1313] = 8'b10110100;
		img[1312] = 8'b10010000;
		img[1311] = 8'b01010010;
		img[1310] = 8'b01110110;
		img[1309] = 8'b10011100;
		img[1308] = 8'b10011010;
		img[1307] = 8'b01101100;
		img[1306] = 8'b01111001;
		img[1305] = 8'b01111100;
		img[1304] = 8'b01110110;
		img[1303] = 8'b00110010;
		img[1302] = 8'b00110100;
		img[1301] = 8'b01100010;
		img[1300] = 8'b00011000;
		img[1299] = 8'b01110001;
		img[1298] = 8'b11001100;
		img[1297] = 8'b01100110;
		img[1296] = 8'b00010000;
		img[1295] = 8'b00000001;
		img[1294] = 8'b00011011;
		img[1293] = 8'b00100001;
		img[1292] = 8'b10001101;
		img[1291] = 8'b01011100;
		img[1290] = 8'b00111100;
		img[1289] = 8'b01000101;
		img[1288] = 8'b00010101;
		img[1287] = 8'b00001011;
		img[1286] = 8'b00011001;
		img[1285] = 8'b00111111;
		img[1284] = 8'b00111101;
		img[1283] = 8'b00100010;
		img[1282] = 8'b00010000;
		img[1281] = 8'b00011101;
		img[1280] = 8'b01001010;
		img[1279] = 8'b00001100;
		img[1278] = 8'b00010001;
		img[1277] = 8'b00100100;
		img[1276] = 8'b00100100;
		img[1275] = 8'b00100101;
		img[1274] = 8'b00001010;
		img[1273] = 8'b00100010;
		img[1272] = 8'b00011101;
		img[1271] = 8'b01000001;
		img[1270] = 8'b01010011;
		img[1269] = 8'b01110111;
		img[1268] = 8'b01101110;
		img[1267] = 8'b01110111;
		img[1266] = 8'b10110001;
		img[1265] = 8'b11010000;
		img[1264] = 8'b11010101;
		img[1263] = 8'b11011110;
		img[1262] = 8'b11011001;
		img[1261] = 8'b11011111;
		img[1260] = 8'b11100000;
		img[1259] = 8'b11001010;
		img[1258] = 8'b11011000;
		img[1257] = 8'b10100111;
		img[1256] = 8'b10110010;
		img[1255] = 8'b01011101;
		img[1254] = 8'b00010111;
		img[1253] = 8'b00000101;
		img[1252] = 8'b00011101;
		img[1251] = 8'b11001001;
		img[1250] = 8'b11011001;
		img[1249] = 8'b10110111;
		img[1248] = 8'b10101001;
		img[1247] = 8'b01010011;
		img[1246] = 8'b01101100;
		img[1245] = 8'b11000110;
		img[1244] = 8'b10010101;
		img[1243] = 8'b01011111;
		img[1242] = 8'b10001110;
		img[1241] = 8'b10010001;
		img[1240] = 8'b01111010;
		img[1239] = 8'b00111000;
		img[1238] = 8'b00111010;
		img[1237] = 8'b01011110;
		img[1236] = 8'b00010101;
		img[1235] = 8'b01111010;
		img[1234] = 8'b10001101;
		img[1233] = 8'b10110111;
		img[1232] = 8'b00111000;
		img[1231] = 8'b00010110;
		img[1230] = 8'b00001101;
		img[1229] = 8'b01000101;
		img[1228] = 8'b10010111;
		img[1227] = 8'b01100111;
		img[1226] = 8'b00000001;
		img[1225] = 8'b11010010;
		img[1224] = 8'b01001110;
		img[1223] = 8'b00100111;
		img[1222] = 8'b00011000;
		img[1221] = 8'b01011000;
		img[1220] = 8'b01001001;
		img[1219] = 8'b00001011;
		img[1218] = 8'b00010111;
		img[1217] = 8'b00111011;
		img[1216] = 8'b00111011;
		img[1215] = 8'b00000111;
		img[1214] = 8'b00000101;
		img[1213] = 8'b00011010;
		img[1212] = 8'b00010110;
		img[1211] = 8'b00011001;
		img[1210] = 8'b00001010;
		img[1209] = 8'b00001111;
		img[1208] = 8'b00011011;
		img[1207] = 8'b00110000;
		img[1206] = 8'b01000011;
		img[1205] = 8'b01100111;
		img[1204] = 8'b01101000;
		img[1203] = 8'b01101010;
		img[1202] = 8'b10110000;
		img[1201] = 8'b11100001;
		img[1200] = 8'b11111001;
		img[1199] = 8'b11101110;
		img[1198] = 8'b11110101;
		img[1197] = 8'b11100011;
		img[1196] = 8'b11011110;
		img[1195] = 8'b11101011;
		img[1194] = 8'b11100111;
		img[1193] = 8'b11010000;
		img[1192] = 8'b10110011;
		img[1191] = 8'b10000011;
		img[1190] = 8'b00100001;
		img[1189] = 8'b00001110;
		img[1188] = 8'b00011000;
		img[1187] = 8'b10111111;
		img[1186] = 8'b11000111;
		img[1185] = 8'b11000001;
		img[1184] = 8'b10111110;
		img[1183] = 8'b01101011;
		img[1182] = 8'b10000110;
		img[1181] = 8'b11011110;
		img[1180] = 8'b10001111;
		img[1179] = 8'b01110110;
		img[1178] = 8'b10001110;
		img[1177] = 8'b10100101;
		img[1176] = 8'b10011000;
		img[1175] = 8'b01010100;
		img[1174] = 8'b00111011;
		img[1173] = 8'b01100100;
		img[1172] = 8'b00000111;
		img[1171] = 8'b11000000;
		img[1170] = 8'b10100100;
		img[1169] = 8'b11011001;
		img[1168] = 8'b01111010;
		img[1167] = 8'b00110000;
		img[1166] = 8'b00010000;
		img[1165] = 8'b00101100;
		img[1164] = 8'b01110011;
		img[1163] = 8'b01100111;
		img[1162] = 8'b01011111;
		img[1161] = 8'b01111101;
		img[1160] = 8'b10010111;
		img[1159] = 8'b10011011;
		img[1158] = 8'b00101000;
		img[1157] = 8'b10010010;
		img[1156] = 8'b10010111;
		img[1155] = 8'b00000000;
		img[1154] = 8'b00001111;
		img[1153] = 8'b00100010;
		img[1152] = 8'b01001010;
		img[1151] = 8'b00010011;
		img[1150] = 8'b00000000;
		img[1149] = 8'b00001011;
		img[1148] = 8'b00000110;
		img[1147] = 8'b00000010;
		img[1146] = 8'b00001011;
		img[1145] = 8'b00001000;
		img[1144] = 8'b00000011;
		img[1143] = 8'b00010101;
		img[1142] = 8'b00111101;
		img[1141] = 8'b01010101;
		img[1140] = 8'b01010110;
		img[1139] = 8'b01100010;
		img[1138] = 8'b10111111;
		img[1137] = 8'b10100010;
		img[1136] = 8'b11001001;
		img[1135] = 8'b11111111;
		img[1134] = 8'b11001111;
		img[1133] = 8'b11111111;
		img[1132] = 8'b11111011;
		img[1131] = 8'b11111101;
		img[1130] = 8'b11100111;
		img[1129] = 8'b11111001;
		img[1128] = 8'b11101101;
		img[1127] = 8'b10111011;
		img[1126] = 8'b01000000;
		img[1125] = 8'b00001101;
		img[1124] = 8'b00011000;
		img[1123] = 8'b10111011;
		img[1122] = 8'b10111100;
		img[1121] = 8'b11010000;
		img[1120] = 8'b11011001;
		img[1119] = 8'b10010111;
		img[1118] = 8'b10101101;
		img[1117] = 8'b11111010;
		img[1116] = 8'b10111110;
		img[1115] = 8'b10101011;
		img[1114] = 8'b11000010;
		img[1113] = 8'b10101101;
		img[1112] = 8'b10111011;
		img[1111] = 8'b01101001;
		img[1110] = 8'b01000101;
		img[1109] = 8'b01101010;
		img[1108] = 8'b00011101;
		img[1107] = 8'b00110010;
		img[1106] = 8'b01111100;
		img[1105] = 8'b10010111;
		img[1104] = 8'b10100010;
		img[1103] = 8'b00011101;
		img[1102] = 8'b01000011;
		img[1101] = 8'b00111101;
		img[1100] = 8'b10011111;
		img[1099] = 8'b01011011;
		img[1098] = 8'b01101111;
		img[1097] = 8'b01110010;
		img[1096] = 8'b01011101;
		img[1095] = 8'b00111000;
		img[1094] = 8'b10011010;
		img[1093] = 8'b10000110;
		img[1092] = 8'b10000110;
		img[1091] = 8'b10001001;
		img[1090] = 8'b00011000;
		img[1089] = 8'b00011100;
		img[1088] = 8'b00111011;
		img[1087] = 8'b00000100;
		img[1086] = 8'b00000000;
		img[1085] = 8'b00001111;
		img[1084] = 8'b00011010;
		img[1083] = 8'b00001001;
		img[1082] = 8'b00000000;
		img[1081] = 8'b00000000;
		img[1080] = 8'b00000010;
		img[1079] = 8'b00010100;
		img[1078] = 8'b00011010;
		img[1077] = 8'b01000000;
		img[1076] = 8'b01010100;
		img[1075] = 8'b10000000;
		img[1074] = 8'b11001110;
		img[1073] = 8'b10100001;
		img[1072] = 8'b10100001;
		img[1071] = 8'b10011010;
		img[1070] = 8'b10101000;
		img[1069] = 8'b10101110;
		img[1068] = 8'b10111111;
		img[1067] = 8'b11000011;
		img[1066] = 8'b10111001;
		img[1065] = 8'b11010111;
		img[1064] = 8'b11110000;
		img[1063] = 8'b11111111;
		img[1062] = 8'b11110000;
		img[1061] = 8'b01000001;
		img[1060] = 8'b00110110;
		img[1059] = 8'b11000101;
		img[1058] = 8'b10111000;
		img[1057] = 8'b11101011;
		img[1056] = 8'b11101000;
		img[1055] = 8'b11101000;
		img[1054] = 8'b11111111;
		img[1053] = 8'b11111111;
		img[1052] = 8'b11111111;
		img[1051] = 8'b11110100;
		img[1050] = 8'b11110110;
		img[1049] = 8'b11111111;
		img[1048] = 8'b11101101;
		img[1047] = 8'b11001100;
		img[1046] = 8'b01010001;
		img[1045] = 8'b01110000;
		img[1044] = 8'b00110101;
		img[1043] = 8'b01101001;
		img[1042] = 8'b10100000;
		img[1041] = 8'b10110110;
		img[1040] = 8'b10010010;
		img[1039] = 8'b01000011;
		img[1038] = 8'b00110110;
		img[1037] = 8'b10010000;
		img[1036] = 8'b11011001;
		img[1035] = 8'b11000100;
		img[1034] = 8'b01100001;
		img[1033] = 8'b01000101;
		img[1032] = 8'b01110000;
		img[1031] = 8'b00011011;
		img[1030] = 8'b11010010;
		img[1029] = 8'b11101111;
		img[1028] = 8'b10001011;
		img[1027] = 8'b10001000;
		img[1026] = 8'b10001011;
		img[1025] = 8'b11010000;
		img[1024] = 8'b01000101;
		img[1023] = 8'b00001101;
		img[1022] = 8'b00001001;
		img[1021] = 8'b00001011;
		img[1020] = 8'b00000000;
		img[1019] = 8'b00000000;
		img[1018] = 8'b00000101;
		img[1017] = 8'b00000000;
		img[1016] = 8'b00001000;
		img[1015] = 8'b00000000;
		img[1014] = 8'b00011100;
		img[1013] = 8'b00101001;
		img[1012] = 8'b10111100;
		img[1011] = 8'b10101101;
		img[1010] = 8'b10100110;
		img[1009] = 8'b10001010;
		img[1008] = 8'b10000111;
		img[1007] = 8'b10000101;
		img[1006] = 8'b10000101;
		img[1005] = 8'b10000011;
		img[1004] = 8'b01101101;
		img[1003] = 8'b01010000;
		img[1002] = 8'b00111001;
		img[1001] = 8'b00101100;
		img[1000] = 8'b00011111;
		img[999] = 8'b00010010;
		img[998] = 8'b00010000;
		img[997] = 8'b00111000;
		img[996] = 8'b00111101;
		img[995] = 8'b00000011;
		img[994] = 8'b00111110;
		img[993] = 8'b00110001;
		img[992] = 8'b00110100;
		img[991] = 8'b00111111;
		img[990] = 8'b01110011;
		img[989] = 8'b01001110;
		img[988] = 8'b01110010;
		img[987] = 8'b01110100;
		img[986] = 8'b01111001;
		img[985] = 8'b01010011;
		img[984] = 8'b01110100;
		img[983] = 8'b01110100;
		img[982] = 8'b10110101;
		img[981] = 8'b10111010;
		img[980] = 8'b00101101;
		img[979] = 8'b01001101;
		img[978] = 8'b00100000;
		img[977] = 8'b01000001;
		img[976] = 8'b11000001;
		img[975] = 8'b01110101;
		img[974] = 8'b00111011;
		img[973] = 8'b01011111;
		img[972] = 8'b00110010;
		img[971] = 8'b01000111;
		img[970] = 8'b10110010;
		img[969] = 8'b01101111;
		img[968] = 8'b00001101;
		img[967] = 8'b00001111;
		img[966] = 8'b00111110;
		img[965] = 8'b01101101;
		img[964] = 8'b00001100;
		img[963] = 8'b01000000;
		img[962] = 8'b00111001;
		img[961] = 8'b00111110;
		img[960] = 8'b10000101;
		img[959] = 8'b00001111;
		img[958] = 8'b00001111;
		img[957] = 8'b00000101;
		img[956] = 8'b00000100;
		img[955] = 8'b00000100;
		img[954] = 8'b00011001;
		img[953] = 8'b00011011;
		img[952] = 8'b00001011;
		img[951] = 8'b00000000;
		img[950] = 8'b00001101;
		img[949] = 8'b00011110;
		img[948] = 8'b10111000;
		img[947] = 8'b10101101;
		img[946] = 8'b10011110;
		img[945] = 8'b10010001;
		img[944] = 8'b10000110;
		img[943] = 8'b10000111;
		img[942] = 8'b10000000;
		img[941] = 8'b01111101;
		img[940] = 8'b01111101;
		img[939] = 8'b01111000;
		img[938] = 8'b01101010;
		img[937] = 8'b01010010;
		img[936] = 8'b00110101;
		img[935] = 8'b00100111;
		img[934] = 8'b00100000;
		img[933] = 8'b00010110;
		img[932] = 8'b00100000;
		img[931] = 8'b00101001;
		img[930] = 8'b00110101;
		img[929] = 8'b01000011;
		img[928] = 8'b01001001;
		img[927] = 8'b01000111;
		img[926] = 8'b00110110;
		img[925] = 8'b00101110;
		img[924] = 8'b00100000;
		img[923] = 8'b00100110;
		img[922] = 8'b00111001;
		img[921] = 8'b01011110;
		img[920] = 8'b01110011;
		img[919] = 8'b01100010;
		img[918] = 8'b01010110;
		img[917] = 8'b01011000;
		img[916] = 8'b10000000;
		img[915] = 8'b01111010;
		img[914] = 8'b10000001;
		img[913] = 8'b00101100;
		img[912] = 8'b01100101;
		img[911] = 8'b00110111;
		img[910] = 8'b00111011;
		img[909] = 8'b00101111;
		img[908] = 8'b00110000;
		img[907] = 8'b01110010;
		img[906] = 8'b01011111;
		img[905] = 8'b10100001;
		img[904] = 8'b10110111;
		img[903] = 8'b00010101;
		img[902] = 8'b11000110;
		img[901] = 8'b10011001;
		img[900] = 8'b01111011;
		img[899] = 8'b01010100;
		img[898] = 8'b01111011;
		img[897] = 8'b01101001;
		img[896] = 8'b00101010;
		img[895] = 8'b00000000;
		img[894] = 8'b00000000;
		img[893] = 8'b00001011;
		img[892] = 8'b00001000;
		img[891] = 8'b00010011;
		img[890] = 8'b00001011;
		img[889] = 8'b00101101;
		img[888] = 8'b00000011;
		img[887] = 8'b00010011;
		img[886] = 8'b00000010;
		img[885] = 8'b00001000;
		img[884] = 8'b01100100;
		img[883] = 8'b10110110;
		img[882] = 8'b10100111;
		img[881] = 8'b10010110;
		img[880] = 8'b10010101;
		img[879] = 8'b10001011;
		img[878] = 8'b10001110;
		img[877] = 8'b10010010;
		img[876] = 8'b10010011;
		img[875] = 8'b10001100;
		img[874] = 8'b10000010;
		img[873] = 8'b01110010;
		img[872] = 8'b01100011;
		img[871] = 8'b01011010;
		img[870] = 8'b01100011;
		img[869] = 8'b01011010;
		img[868] = 8'b01011011;
		img[867] = 8'b01101000;
		img[866] = 8'b01101110;
		img[865] = 8'b01110010;
		img[864] = 8'b01100100;
		img[863] = 8'b01010000;
		img[862] = 8'b01000111;
		img[861] = 8'b00110101;
		img[860] = 8'b00011011;
		img[859] = 8'b00001111;
		img[858] = 8'b00011011;
		img[857] = 8'b00101111;
		img[856] = 8'b01001110;
		img[855] = 8'b01011101;
		img[854] = 8'b01100001;
		img[853] = 8'b01100000;
		img[852] = 8'b01011110;
		img[851] = 8'b01100111;
		img[850] = 8'b01111111;
		img[849] = 8'b01011011;
		img[848] = 8'b00010101;
		img[847] = 8'b00100001;
		img[846] = 8'b01001101;
		img[845] = 8'b00010100;
		img[844] = 8'b01010111;
		img[843] = 8'b01010101;
		img[842] = 8'b01010111;
		img[841] = 8'b01100011;
		img[840] = 8'b10000111;
		img[839] = 8'b10110011;
		img[838] = 8'b11001010;
		img[837] = 8'b11001000;
		img[836] = 8'b10010101;
		img[835] = 8'b01001100;
		img[834] = 8'b11010101;
		img[833] = 8'b01110001;
		img[832] = 8'b10010010;
		img[831] = 8'b00010010;
		img[830] = 8'b00010011;
		img[829] = 8'b00001010;
		img[828] = 8'b00010001;
		img[827] = 8'b00001011;
		img[826] = 8'b00000101;
		img[825] = 8'b00011101;
		img[824] = 8'b00000100;
		img[823] = 8'b00001100;
		img[822] = 8'b01011011;
		img[821] = 8'b10001001;
		img[820] = 8'b10111001;
		img[819] = 8'b11001111;
		img[818] = 8'b10111110;
		img[817] = 8'b10111001;
		img[816] = 8'b10111101;
		img[815] = 8'b10111010;
		img[814] = 8'b10111010;
		img[813] = 8'b10111000;
		img[812] = 8'b10110111;
		img[811] = 8'b10101010;
		img[810] = 8'b10100011;
		img[809] = 8'b10010111;
		img[808] = 8'b10010011;
		img[807] = 8'b10001011;
		img[806] = 8'b10000111;
		img[805] = 8'b10001001;
		img[804] = 8'b10001001;
		img[803] = 8'b01111111;
		img[802] = 8'b10000010;
		img[801] = 8'b01111001;
		img[800] = 8'b01110001;
		img[799] = 8'b01100101;
		img[798] = 8'b01100001;
		img[797] = 8'b01010010;
		img[796] = 8'b01001000;
		img[795] = 8'b01001010;
		img[794] = 8'b01010010;
		img[793] = 8'b01100111;
		img[792] = 8'b01110110;
		img[791] = 8'b10000100;
		img[790] = 8'b01111000;
		img[789] = 8'b01101111;
		img[788] = 8'b01101010;
		img[787] = 8'b01110010;
		img[786] = 8'b01110010;
		img[785] = 8'b01001010;
		img[784] = 8'b01000001;
		img[783] = 8'b01000111;
		img[782] = 8'b10000010;
		img[781] = 8'b00101110;
		img[780] = 8'b00110101;
		img[779] = 8'b01101110;
		img[778] = 8'b01111111;
		img[777] = 8'b01111100;
		img[776] = 8'b10000000;
		img[775] = 8'b10001111;
		img[774] = 8'b10011010;
		img[773] = 8'b11000001;
		img[772] = 8'b10001011;
		img[771] = 8'b01001110;
		img[770] = 8'b10100001;
		img[769] = 8'b01010100;
		img[768] = 8'b10111111;
		img[767] = 8'b00000100;
		img[766] = 8'b00000111;
		img[765] = 8'b00001000;
		img[764] = 8'b00001010;
		img[763] = 8'b00011001;
		img[762] = 8'b00000000;
		img[761] = 8'b00000000;
		img[760] = 8'b00000111;
		img[759] = 8'b00100001;
		img[758] = 8'b11010111;
		img[757] = 8'b11101101;
		img[756] = 8'b11101000;
		img[755] = 8'b11011111;
		img[754] = 8'b11010111;
		img[753] = 8'b11011011;
		img[752] = 8'b11011100;
		img[751] = 8'b11100001;
		img[750] = 8'b11100100;
		img[749] = 8'b11100000;
		img[748] = 8'b11011000;
		img[747] = 8'b11000101;
		img[746] = 8'b10111010;
		img[745] = 8'b10110011;
		img[744] = 8'b10110110;
		img[743] = 8'b10110101;
		img[742] = 8'b10110011;
		img[741] = 8'b10110000;
		img[740] = 8'b10110010;
		img[739] = 8'b10111000;
		img[738] = 8'b10101000;
		img[737] = 8'b10100101;
		img[736] = 8'b10011101;
		img[735] = 8'b10011101;
		img[734] = 8'b10011001;
		img[733] = 8'b10011000;
		img[732] = 8'b10010011;
		img[731] = 8'b10010101;
		img[730] = 8'b10010010;
		img[729] = 8'b10011111;
		img[728] = 8'b10011011;
		img[727] = 8'b10011101;
		img[726] = 8'b10100111;
		img[725] = 8'b10101001;
		img[724] = 8'b10101100;
		img[723] = 8'b10101010;
		img[722] = 8'b10110010;
		img[721] = 8'b11000111;
		img[720] = 8'b11000010;
		img[719] = 8'b10110110;
		img[718] = 8'b10110011;
		img[717] = 8'b10010000;
		img[716] = 8'b00000000;
		img[715] = 8'b01000001;
		img[714] = 8'b10000110;
		img[713] = 8'b10011110;
		img[712] = 8'b10100101;
		img[711] = 8'b10110010;
		img[710] = 8'b10111001;
		img[709] = 8'b11001010;
		img[708] = 8'b11000010;
		img[707] = 8'b00100000;
		img[706] = 8'b11001110;
		img[705] = 8'b10100100;
		img[704] = 8'b00100101;
		img[703] = 8'b00001001;
		img[702] = 8'b00010011;
		img[701] = 8'b00001010;
		img[700] = 8'b00000000;
		img[699] = 8'b00001011;
		img[698] = 8'b00000000;
		img[697] = 8'b00000100;
		img[696] = 8'b00001000;
		img[695] = 8'b00101001;
		img[694] = 8'b01110110;
		img[693] = 8'b11100110;
		img[692] = 8'b11100010;
		img[691] = 8'b11011011;
		img[690] = 8'b11100101;
		img[689] = 8'b11100100;
		img[688] = 8'b11101011;
		img[687] = 8'b11101111;
		img[686] = 8'b11101101;
		img[685] = 8'b11100001;
		img[684] = 8'b11010110;
		img[683] = 8'b11001000;
		img[682] = 8'b10111110;
		img[681] = 8'b10110111;
		img[680] = 8'b10110111;
		img[679] = 8'b10111110;
		img[678] = 8'b11001111;
		img[677] = 8'b11010110;
		img[676] = 8'b11010010;
		img[675] = 8'b11010111;
		img[674] = 8'b11001101;
		img[673] = 8'b11001011;
		img[672] = 8'b11000010;
		img[671] = 8'b11000111;
		img[670] = 8'b11010000;
		img[669] = 8'b11010001;
		img[668] = 8'b11010011;
		img[667] = 8'b11010001;
		img[666] = 8'b11001100;
		img[665] = 8'b10111000;
		img[664] = 8'b10111011;
		img[663] = 8'b10101111;
		img[662] = 8'b10111001;
		img[661] = 8'b10110111;
		img[660] = 8'b10111111;
		img[659] = 8'b11001000;
		img[658] = 8'b11010000;
		img[657] = 8'b11011010;
		img[656] = 8'b11010111;
		img[655] = 8'b11010110;
		img[654] = 8'b11001100;
		img[653] = 8'b11010010;
		img[652] = 8'b01010100;
		img[651] = 8'b01011010;
		img[650] = 8'b10011101;
		img[649] = 8'b11000110;
		img[648] = 8'b11000111;
		img[647] = 8'b11010010;
		img[646] = 8'b11001011;
		img[645] = 8'b11010011;
		img[644] = 8'b11011101;
		img[643] = 8'b11101011;
		img[642] = 8'b11100001;
		img[641] = 8'b11110100;
		img[640] = 8'b10101001;
		img[639] = 8'b00000000;
		img[638] = 8'b00010010;
		img[637] = 8'b00001001;
		img[636] = 8'b00100111;
		img[635] = 8'b00000100;
		img[634] = 8'b00010011;
		img[633] = 8'b00000000;
		img[632] = 8'b00101010;
		img[631] = 8'b00000100;
		img[630] = 8'b00101001;
		img[629] = 8'b10100111;
		img[628] = 8'b10101001;
		img[627] = 8'b10110001;
		img[626] = 8'b10111110;
		img[625] = 8'b11000001;
		img[624] = 8'b11000111;
		img[623] = 8'b11001101;
		img[622] = 8'b11001110;
		img[621] = 8'b11000100;
		img[620] = 8'b10110010;
		img[619] = 8'b10100111;
		img[618] = 8'b10011101;
		img[617] = 8'b10011111;
		img[616] = 8'b10100111;
		img[615] = 8'b10101110;
		img[614] = 8'b10110011;
		img[613] = 8'b11000101;
		img[612] = 8'b11001001;
		img[611] = 8'b11000001;
		img[610] = 8'b11000101;
		img[609] = 8'b11001001;
		img[608] = 8'b11010110;
		img[607] = 8'b11101100;
		img[606] = 8'b11101111;
		img[605] = 8'b11110010;
		img[604] = 8'b11101100;
		img[603] = 8'b11101000;
		img[602] = 8'b11010010;
		img[601] = 8'b11000010;
		img[600] = 8'b10111100;
		img[599] = 8'b10111101;
		img[598] = 8'b11000101;
		img[597] = 8'b11001111;
		img[596] = 8'b11011101;
		img[595] = 8'b11011110;
		img[594] = 8'b11100100;
		img[593] = 8'b11011011;
		img[592] = 8'b11011001;
		img[591] = 8'b11011101;
		img[590] = 8'b11010011;
		img[589] = 8'b11101011;
		img[588] = 8'b01110001;
		img[587] = 8'b10111110;
		img[586] = 8'b11101001;
		img[585] = 8'b11100101;
		img[584] = 8'b11101011;
		img[583] = 8'b11101100;
		img[582] = 8'b11110100;
		img[581] = 8'b11110001;
		img[580] = 8'b11110000;
		img[579] = 8'b11101101;
		img[578] = 8'b11110000;
		img[577] = 8'b11110110;
		img[576] = 8'b11110100;
		img[575] = 8'b01001001;
		img[574] = 8'b01101101;
		img[573] = 8'b00000000;
		img[572] = 8'b00000000;
		img[571] = 8'b00000100;
		img[570] = 8'b00000000;
		img[569] = 8'b00001001;
		img[568] = 8'b00000000;
		img[567] = 8'b00001001;
		img[566] = 8'b00000001;
		img[565] = 8'b10010111;
		img[564] = 8'b10100111;
		img[563] = 8'b10101110;
		img[562] = 8'b10110101;
		img[561] = 8'b10111000;
		img[560] = 8'b10111000;
		img[559] = 8'b10111010;
		img[558] = 8'b10110000;
		img[557] = 8'b10011111;
		img[556] = 8'b10010000;
		img[555] = 8'b10010111;
		img[554] = 8'b10011000;
		img[553] = 8'b10010100;
		img[552] = 8'b10001111;
		img[551] = 8'b10000110;
		img[550] = 8'b10000011;
		img[549] = 8'b10001011;
		img[548] = 8'b10001110;
		img[547] = 8'b10001000;
		img[546] = 8'b01111010;
		img[545] = 8'b01110101;
		img[544] = 8'b01111011;
		img[543] = 8'b10011000;
		img[542] = 8'b11000111;
		img[541] = 8'b11011000;
		img[540] = 8'b11011101;
		img[539] = 8'b11001011;
		img[538] = 8'b10010110;
		img[537] = 8'b10000100;
		img[536] = 8'b10000110;
		img[535] = 8'b10011000;
		img[534] = 8'b10110111;
		img[533] = 8'b11001111;
		img[532] = 8'b11011110;
		img[531] = 8'b11101100;
		img[530] = 8'b11101000;
		img[529] = 8'b11100001;
		img[528] = 8'b11011011;
		img[527] = 8'b11100011;
		img[526] = 8'b11101011;
		img[525] = 8'b11101110;
		img[524] = 8'b11001111;
		img[523] = 8'b11110011;
		img[522] = 8'b11101110;
		img[521] = 8'b11101111;
		img[520] = 8'b11110110;
		img[519] = 8'b11110111;
		img[518] = 8'b11111000;
		img[517] = 8'b11110111;
		img[516] = 8'b11111000;
		img[515] = 8'b11111010;
		img[514] = 8'b11111110;
		img[513] = 8'b11111001;
		img[512] = 8'b11111110;
		img[511] = 8'b10110011;
		img[510] = 8'b00111101;
		img[509] = 8'b00110011;
		img[508] = 8'b00110010;
		img[507] = 8'b00000110;
		img[506] = 8'b00000000;
		img[505] = 8'b00000000;
		img[504] = 8'b00000011;
		img[503] = 8'b00000011;
		img[502] = 8'b01100000;
		img[501] = 8'b10111010;
		img[500] = 8'b11000110;
		img[499] = 8'b11000111;
		img[498] = 8'b11000010;
		img[497] = 8'b10111000;
		img[496] = 8'b10101011;
		img[495] = 8'b10110010;
		img[494] = 8'b10101100;
		img[493] = 8'b10100010;
		img[492] = 8'b10010101;
		img[491] = 8'b10001010;
		img[490] = 8'b10000010;
		img[489] = 8'b01101111;
		img[488] = 8'b01010110;
		img[487] = 8'b00110000;
		img[486] = 8'b00100000;
		img[485] = 8'b00100000;
		img[484] = 8'b00101111;
		img[483] = 8'b01001010;
		img[482] = 8'b01101000;
		img[481] = 8'b01110011;
		img[480] = 8'b01111000;
		img[479] = 8'b01101111;
		img[478] = 8'b01101010;
		img[477] = 8'b01101101;
		img[476] = 8'b01110110;
		img[475] = 8'b10000000;
		img[474] = 8'b10000110;
		img[473] = 8'b10001100;
		img[472] = 8'b10010111;
		img[471] = 8'b10101011;
		img[470] = 8'b11000011;
		img[469] = 8'b11011001;
		img[468] = 8'b11100101;
		img[467] = 8'b11101011;
		img[466] = 8'b11101100;
		img[465] = 8'b11101011;
		img[464] = 8'b11101100;
		img[463] = 8'b11110010;
		img[462] = 8'b11110011;
		img[461] = 8'b11110100;
		img[460] = 8'b11111011;
		img[459] = 8'b11110101;
		img[458] = 8'b11110100;
		img[457] = 8'b11110001;
		img[456] = 8'b11110011;
		img[455] = 8'b11110011;
		img[454] = 8'b11110111;
		img[453] = 8'b11111001;
		img[452] = 8'b11111011;
		img[451] = 8'b11111101;
		img[450] = 8'b11111111;
		img[449] = 8'b11111110;
		img[448] = 8'b11111100;
		img[447] = 8'b11011101;
		img[446] = 8'b11001111;
		img[445] = 8'b10010101;
		img[444] = 8'b10101100;
		img[443] = 8'b10001000;
		img[442] = 8'b00001100;
		img[441] = 8'b00110100;
		img[440] = 8'b00100000;
		img[439] = 8'b00010100;
		img[438] = 8'b10111110;
		img[437] = 8'b11000010;
		img[436] = 8'b10111111;
		img[435] = 8'b11000010;
		img[434] = 8'b10111111;
		img[433] = 8'b10111110;
		img[432] = 8'b10111001;
		img[431] = 8'b10111110;
		img[430] = 8'b10111100;
		img[429] = 8'b10110010;
		img[428] = 8'b10010100;
		img[427] = 8'b01101101;
		img[426] = 8'b01010000;
		img[425] = 8'b01000011;
		img[424] = 8'b00111100;
		img[423] = 8'b00100110;
		img[422] = 8'b00001110;
		img[421] = 8'b00000010;
		img[420] = 8'b00000010;
		img[419] = 8'b00010100;
		img[418] = 8'b00110110;
		img[417] = 8'b01010100;
		img[416] = 8'b01100111;
		img[415] = 8'b01101000;
		img[414] = 8'b01101111;
		img[413] = 8'b01111110;
		img[412] = 8'b10001100;
		img[411] = 8'b10010101;
		img[410] = 8'b10011111;
		img[409] = 8'b10101111;
		img[408] = 8'b11000000;
		img[407] = 8'b11000110;
		img[406] = 8'b11001011;
		img[405] = 8'b11010001;
		img[404] = 8'b11011001;
		img[403] = 8'b11100001;
		img[402] = 8'b11100100;
		img[401] = 8'b11101011;
		img[400] = 8'b11110101;
		img[399] = 8'b11110101;
		img[398] = 8'b11111000;
		img[397] = 8'b11111011;
		img[396] = 8'b11111011;
		img[395] = 8'b11111100;
		img[394] = 8'b11111100;
		img[393] = 8'b11111001;
		img[392] = 8'b11110010;
		img[391] = 8'b11110101;
		img[390] = 8'b11110011;
		img[389] = 8'b11110011;
		img[388] = 8'b11110111;
		img[387] = 8'b11111001;
		img[386] = 8'b11110011;
		img[385] = 8'b11101101;
		img[384] = 8'b11101010;
		img[383] = 8'b11011100;
		img[382] = 8'b11011110;
		img[381] = 8'b11010100;
		img[380] = 8'b11010100;
		img[379] = 8'b10101101;
		img[378] = 8'b01110110;
		img[377] = 8'b11001100;
		img[376] = 8'b11010100;
		img[375] = 8'b10111100;
		img[374] = 8'b11001001;
		img[373] = 8'b11000011;
		img[372] = 8'b11010000;
		img[371] = 8'b11001010;
		img[370] = 8'b11000100;
		img[369] = 8'b10111100;
		img[368] = 8'b10111110;
		img[367] = 8'b11000010;
		img[366] = 8'b10110101;
		img[365] = 8'b10100010;
		img[364] = 8'b10001000;
		img[363] = 8'b01101010;
		img[362] = 8'b01010011;
		img[361] = 8'b01000011;
		img[360] = 8'b00111000;
		img[359] = 8'b00101001;
		img[358] = 8'b00010110;
		img[357] = 8'b00001110;
		img[356] = 8'b00010011;
		img[355] = 8'b00101001;
		img[354] = 8'b01001010;
		img[353] = 8'b01100011;
		img[352] = 8'b01110100;
		img[351] = 8'b01101100;
		img[350] = 8'b01011111;
		img[349] = 8'b01011001;
		img[348] = 8'b01100110;
		img[347] = 8'b01111111;
		img[346] = 8'b10010101;
		img[345] = 8'b10011011;
		img[344] = 8'b10011011;
		img[343] = 8'b10011000;
		img[342] = 8'b10010101;
		img[341] = 8'b10010101;
		img[340] = 8'b10100100;
		img[339] = 8'b10110111;
		img[338] = 8'b11001000;
		img[337] = 8'b11011001;
		img[336] = 8'b11101010;
		img[335] = 8'b11110010;
		img[334] = 8'b11110101;
		img[333] = 8'b11111101;
		img[332] = 8'b11111011;
		img[331] = 8'b11111100;
		img[330] = 8'b11110111;
		img[329] = 8'b11111001;
		img[328] = 8'b11111001;
		img[327] = 8'b11111100;
		img[326] = 8'b11111101;
		img[325] = 8'b11110110;
		img[324] = 8'b11011100;
		img[323] = 8'b10101110;
		img[322] = 8'b10000111;
		img[321] = 8'b10000100;
		img[320] = 8'b10010101;
		img[319] = 8'b11101001;
		img[318] = 8'b11100101;
		img[317] = 8'b11011111;
		img[316] = 8'b11010111;
		img[315] = 8'b11101001;
		img[314] = 8'b11101011;
		img[313] = 8'b11100100;
		img[312] = 8'b11011110;
		img[311] = 8'b11010010;
		img[310] = 8'b11010100;
		img[309] = 8'b11010111;
		img[308] = 8'b11011101;
		img[307] = 8'b11100011;
		img[306] = 8'b11010110;
		img[305] = 8'b11011000;
		img[304] = 8'b11010000;
		img[303] = 8'b11001011;
		img[302] = 8'b10111101;
		img[301] = 8'b10100110;
		img[300] = 8'b10001110;
		img[299] = 8'b01111011;
		img[298] = 8'b01110001;
		img[297] = 8'b01100101;
		img[296] = 8'b01011011;
		img[295] = 8'b01010101;
		img[294] = 8'b01001010;
		img[293] = 8'b01000101;
		img[292] = 8'b01000010;
		img[291] = 8'b01001010;
		img[290] = 8'b01011101;
		img[289] = 8'b01110100;
		img[288] = 8'b10000101;
		img[287] = 8'b10011000;
		img[286] = 8'b10010011;
		img[285] = 8'b10000110;
		img[284] = 8'b01110111;
		img[283] = 8'b01101100;
		img[282] = 8'b01101110;
		img[281] = 8'b01111001;
		img[280] = 8'b10000011;
		img[279] = 8'b10001000;
		img[278] = 8'b10001101;
		img[277] = 8'b10010100;
		img[276] = 8'b10100001;
		img[275] = 8'b10110111;
		img[274] = 8'b11001100;
		img[273] = 8'b11011011;
		img[272] = 8'b11100100;
		img[271] = 8'b11100001;
		img[270] = 8'b11011010;
		img[269] = 8'b11011001;
		img[268] = 8'b11011011;
		img[267] = 8'b11101001;
		img[266] = 8'b11101100;
		img[265] = 8'b11100111;
		img[264] = 8'b11100000;
		img[263] = 8'b11010111;
		img[262] = 8'b11001010;
		img[261] = 8'b10111011;
		img[260] = 8'b10101100;
		img[259] = 8'b10010001;
		img[258] = 8'b01110000;
		img[257] = 8'b01011011;
		img[256] = 8'b01010110;
		img[255] = 8'b11100000;
		img[254] = 8'b11100110;
		img[253] = 8'b11100010;
		img[252] = 8'b11011110;
		img[251] = 8'b11011101;
		img[250] = 8'b11011110;
		img[249] = 8'b11011011;
		img[248] = 8'b11011111;
		img[247] = 8'b11011011;
		img[246] = 8'b11011001;
		img[245] = 8'b11011111;
		img[244] = 8'b11100000;
		img[243] = 8'b11100100;
		img[242] = 8'b11100010;
		img[241] = 8'b11011101;
		img[240] = 8'b11011000;
		img[239] = 8'b11000101;
		img[238] = 8'b10111100;
		img[237] = 8'b10101100;
		img[236] = 8'b10010111;
		img[235] = 8'b10000110;
		img[234] = 8'b01111110;
		img[233] = 8'b01111110;
		img[232] = 8'b01111100;
		img[231] = 8'b01111011;
		img[230] = 8'b01110111;
		img[229] = 8'b01110100;
		img[228] = 8'b01101100;
		img[227] = 8'b01100010;
		img[226] = 8'b01100000;
		img[225] = 8'b01011110;
		img[224] = 8'b01100001;
		img[223] = 8'b10000111;
		img[222] = 8'b10001101;
		img[221] = 8'b10001110;
		img[220] = 8'b10000110;
		img[219] = 8'b01111100;
		img[218] = 8'b01110111;
		img[217] = 8'b01110111;
		img[216] = 8'b01111001;
		img[215] = 8'b10001110;
		img[214] = 8'b10100001;
		img[213] = 8'b10110011;
		img[212] = 8'b11000101;
		img[211] = 8'b11011100;
		img[210] = 8'b11101100;
		img[209] = 8'b11110011;
		img[208] = 8'b11110100;
		img[207] = 8'b11101111;
		img[206] = 8'b11101101;
		img[205] = 8'b11001100;
		img[204] = 8'b10011101;
		img[203] = 8'b10001100;
		img[202] = 8'b10100100;
		img[201] = 8'b10111001;
		img[200] = 8'b11000100;
		img[199] = 8'b10111100;
		img[198] = 8'b10110000;
		img[197] = 8'b10100100;
		img[196] = 8'b10100000;
		img[195] = 8'b10011001;
		img[194] = 8'b10010010;
		img[193] = 8'b10010001;
		img[192] = 8'b10010100;
		img[191] = 8'b11100110;
		img[190] = 8'b11100001;
		img[189] = 8'b11100101;
		img[188] = 8'b11100000;
		img[187] = 8'b11011101;
		img[186] = 8'b11011110;
		img[185] = 8'b11011100;
		img[184] = 8'b11100010;
		img[183] = 8'b11011110;
		img[182] = 8'b11011111;
		img[181] = 8'b11011111;
		img[180] = 8'b11011010;
		img[179] = 8'b11010111;
		img[178] = 8'b11010010;
		img[177] = 8'b11001110;
		img[176] = 8'b11000100;
		img[175] = 8'b10111010;
		img[174] = 8'b10110101;
		img[173] = 8'b10110001;
		img[172] = 8'b10101111;
		img[171] = 8'b10101011;
		img[170] = 8'b10100100;
		img[169] = 8'b10011111;
		img[168] = 8'b10011100;
		img[167] = 8'b10010101;
		img[166] = 8'b10001011;
		img[165] = 8'b10000100;
		img[164] = 8'b01111011;
		img[163] = 8'b01110000;
		img[162] = 8'b01101001;
		img[161] = 8'b01100000;
		img[160] = 8'b01011011;
		img[159] = 8'b01101011;
		img[158] = 8'b01110000;
		img[157] = 8'b01110100;
		img[156] = 8'b01110110;
		img[155] = 8'b01111000;
		img[154] = 8'b01111100;
		img[153] = 8'b10000000;
		img[152] = 8'b10000011;
		img[151] = 8'b10010111;
		img[150] = 8'b10101011;
		img[149] = 8'b11000010;
		img[148] = 8'b11010101;
		img[147] = 8'b11100100;
		img[146] = 8'b11101100;
		img[145] = 8'b11101011;
		img[144] = 8'b11101011;
		img[143] = 8'b11110010;
		img[142] = 8'b11100011;
		img[141] = 8'b11000111;
		img[140] = 8'b10101111;
		img[139] = 8'b10001111;
		img[138] = 8'b01111001;
		img[137] = 8'b01110010;
		img[136] = 8'b10000100;
		img[135] = 8'b10010001;
		img[134] = 8'b10010101;
		img[133] = 8'b10011010;
		img[132] = 8'b10100000;
		img[131] = 8'b10100010;
		img[130] = 8'b10100110;
		img[129] = 8'b10101010;
		img[128] = 8'b10101111;
		img[127] = 8'b11101010;
		img[126] = 8'b11101001;
		img[125] = 8'b11101101;
		img[124] = 8'b11101010;
		img[123] = 8'b11101001;
		img[122] = 8'b11100111;
		img[121] = 8'b11100011;
		img[120] = 8'b11011011;
		img[119] = 8'b11011110;
		img[118] = 8'b11010101;
		img[117] = 8'b11010001;
		img[116] = 8'b10111101;
		img[115] = 8'b10110111;
		img[114] = 8'b10110011;
		img[113] = 8'b10111001;
		img[112] = 8'b10110011;
		img[111] = 8'b10110111;
		img[110] = 8'b10111010;
		img[109] = 8'b11000011;
		img[108] = 8'b11001010;
		img[107] = 8'b11000100;
		img[106] = 8'b10111010;
		img[105] = 8'b10101011;
		img[104] = 8'b10011110;
		img[103] = 8'b10010000;
		img[102] = 8'b10001011;
		img[101] = 8'b10001101;
		img[100] = 8'b10001000;
		img[99] = 8'b10000000;
		img[98] = 8'b01111001;
		img[97] = 8'b01110001;
		img[96] = 8'b01110000;
		img[95] = 8'b01111010;
		img[94] = 8'b10000101;
		img[93] = 8'b10010001;
		img[92] = 8'b10011010;
		img[91] = 8'b10100000;
		img[90] = 8'b10100100;
		img[89] = 8'b10100100;
		img[88] = 8'b10100110;
		img[87] = 8'b10100111;
		img[86] = 8'b10111000;
		img[85] = 8'b11001000;
		img[84] = 8'b11011000;
		img[83] = 8'b11100100;
		img[82] = 8'b11100111;
		img[81] = 8'b11100101;
		img[80] = 8'b11100111;
		img[79] = 8'b11100111;
		img[78] = 8'b11100110;
		img[77] = 8'b11011010;
		img[76] = 8'b11001010;
		img[75] = 8'b10111001;
		img[74] = 8'b10100011;
		img[73] = 8'b10010000;
		img[72] = 8'b10001100;
		img[71] = 8'b10001011;
		img[70] = 8'b10010011;
		img[69] = 8'b10011110;
		img[68] = 8'b10100110;
		img[67] = 8'b10101011;
		img[66] = 8'b10101101;
		img[65] = 8'b10101011;
		img[64] = 8'b10101010;
		img[63] = 8'b11101110;
		img[62] = 8'b11110110;
		img[61] = 8'b11111010;
		img[60] = 8'b11111111;
		img[59] = 8'b11111101;
		img[58] = 8'b11110110;
		img[57] = 8'b11101011;
		img[56] = 8'b11101010;
		img[55] = 8'b11011011;
		img[54] = 8'b11001111;
		img[53] = 8'b10110110;
		img[52] = 8'b10100110;
		img[51] = 8'b10100111;
		img[50] = 8'b10100101;
		img[49] = 8'b10101010;
		img[48] = 8'b10111000;
		img[47] = 8'b11000000;
		img[46] = 8'b11001000;
		img[45] = 8'b11001111;
		img[44] = 8'b11001110;
		img[43] = 8'b11001000;
		img[42] = 8'b10111011;
		img[41] = 8'b10100100;
		img[40] = 8'b10001010;
		img[39] = 8'b10000000;
		img[38] = 8'b01111011;
		img[37] = 8'b10000010;
		img[36] = 8'b10000111;
		img[35] = 8'b10001001;
		img[34] = 8'b10000110;
		img[33] = 8'b01111100;
		img[32] = 8'b01110101;
		img[31] = 8'b01111100;
		img[30] = 8'b10000011;
		img[29] = 8'b10010000;
		img[28] = 8'b10011100;
		img[27] = 8'b10100111;
		img[26] = 8'b10101111;
		img[25] = 8'b10110001;
		img[24] = 8'b10110010;
		img[23] = 8'b10110010;
		img[22] = 8'b10111011;
		img[21] = 8'b11000110;
		img[20] = 8'b11001110;
		img[19] = 8'b11010111;
		img[18] = 8'b11011100;
		img[17] = 8'b11011011;
		img[16] = 8'b11011011;
		img[15] = 8'b11100110;
		img[14] = 8'b11100101;
		img[13] = 8'b11100000;
		img[12] = 8'b11010110;
		img[11] = 8'b11010010;
		img[10] = 8'b10111111;
		img[9] = 8'b10110001;
		img[8] = 8'b10101110;
		img[7] = 8'b10101110;
		img[6] = 8'b10110000;
		img[5] = 8'b10110010;
		img[4] = 8'b10110100;
		img[3] = 8'b10110101;
		img[2] = 8'b10110101;
		img[1] = 8'b10110110;
		img[0] = 8'b10111000;
		

  for(ii=0; ii<120; ii=ii+1) begin
    img[4093-ii][0] <= message[119-ii];
	end
end


reg	[27:0]	counter;
initial	counter = 28'hffffff0;
always @(posedge i_clk)
	counter <= counter + 1'b1;

wire		tx_break, tx_busy;
reg		tx_stb;
reg	[3:0]	tx_index;
reg	[7:0]	tx_data;

assign	tx_break = 1'b0;

initial	tx_index = 12'h0;
always @(posedge i_clk)
	if ((tx_stb)&&(!tx_busy))
		tx_index <= tx_index + 1'b1;
always @(posedge i_clk)
	tx_data <= message[tx_index];

initial	tx_stb = 1'b0;
always @(posedge i_clk)
	if (&counter)
		tx_stb <= 1'b1;
	else if ((tx_stb)&&(!tx_busy)&&(tx_index==4'hf))
		tx_stb <= 1'b0;

// 868 is 115200 Baud, based upon a 100MHz clock
txuartlite #(.TIMING_BITS(10), .CLOCKS_PER_BAUD(868))
	transmitter(i_clk, tx_stb, tx_data, o_uart_tx, tx_busy);

endmodule
////////////////////////////////////////////////////////////////////////////////
//
// Filename: 	txuartlite.v
//
// Project:	wbuart32, a full featured UART with simulator
//
// Purpose:	Transmit outputs over a single UART line.  This particular UART
//		implementation has been extremely simplified: it does not handle
//	generating break conditions, nor does it handle anything other than the
//	8N1 (8 data bits, no parity, 1 stop bit) UART sub-protocol.
//
//	To interface with this module, connect it to your system clock, and
//	pass it the byte of data you wish to transmit.  Strobe the i_wr line
//	high for one cycle, and your data will be off.  Wait until the 'o_busy'
//	line is low before strobing the i_wr line again--this implementation
//	has NO BUFFER, so strobing i_wr while the core is busy will just
//	get ignored.  The output will be placed on the o_txuart output line.
//
//	(I often set both data and strobe on the same clock, and then just leave
//	them set until the busy line is low.  Then I move on to the next piece
//	of data.)
//
// Creator:	Dan Gisselquist, Ph.D.
//		Gisselquist Technology, LLC
//
////////////////////////////////////////////////////////////////////////////////
//
// Copyright (C) 2015-2017, Gisselquist Technology, LLC
//
// This program is free software (firmware): you can redistribute it and/or
// modify it under the terms of  the GNU General Public License as published
// by the Free Software Foundation, either version 3 of the License, or (at
// your option) any later version.
//
// This program is distributed in the hope that it will be useful, but WITHOUT
// ANY WARRANTY; without even the implied warranty of MERCHANTIBILITY or
// FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
// for more details.
//
// You should have received a copy of the GNU General Public License along
// with this program.  (It's in the $(ROOT)/doc directory.  Run make with no
// target there if the PDF file isn't present.)  If not, see
// <http://www.gnu.org/licenses/> for a copy.
//
// License:	GPL, v3, as defined and found on www.gnu.org,
//		http://www.gnu.org/licenses/gpl.html
//
//
////////////////////////////////////////////////////////////////////////////////
//
//
`default_nettype	none
//
`define	TXUL_BIT_ZERO	4'h0
`define	TXUL_BIT_ONE	4'h1
`define	TXUL_BIT_TWO	4'h2
`define	TXUL_BIT_THREE	4'h3
`define	TXUL_BIT_FOUR	4'h4
`define	TXUL_BIT_FIVE	4'h5
`define	TXUL_BIT_SIX	4'h6
`define	TXUL_BIT_SEVEN	4'h7
`define	TXUL_STOP	4'h8
`define	TXUL_IDLE	4'hf
//
//
module txuartlite(i_clk, i_wr, i_data, o_uart_tx, o_busy);
parameter	[4:0]	TIMING_BITS = 5'd24;
localparam		TB = TIMING_BITS;
parameter	[(TB-1):0]	CLOCKS_PER_BAUD = 8; // 24'd868;
parameter	[0:0]	F_OPT_CLK2FFLOGIC = 1'b0;
input	wire		i_clk;
input	wire		i_wr;
input	wire	[7:0]	i_data;
// And the UART input line itself
output	reg		o_uart_tx;
// A line to tell others when we are ready to accept data.  If
// (i_wr)&&(!o_busy) is ever true, then the core has accepted a byte
// for transmission.
output	wire		o_busy;

reg	[(TB-1):0]	baud_counter;
reg	[3:0]	state;
reg	[7:0]	lcl_data;
reg		r_busy, zero_baud_counter;

initial	r_busy = 1'b1;
initial	state  = `TXUL_IDLE;
always @(posedge i_clk)
begin
	if (!zero_baud_counter)
		// r_busy needs to be set coming into here
		r_busy <= 1'b1;
	else if (state > `TXUL_STOP)	// STATE_IDLE
	begin
		state <= `TXUL_IDLE;
		r_busy <= 1'b0;
		if ((i_wr)&&(!r_busy))
		begin	// Immediately start us off with a start bit
			r_busy <= 1'b1;
			state <= `TXUL_BIT_ZERO;
		end
	end else begin
		// One clock tick in each of these states ...
		r_busy <= 1'b1;
		if (state <=`TXUL_STOP) // start bit, 8-d bits, stop-b
			state <= state + 1'b1;
		else
			state <= `TXUL_IDLE;
	end
end

// o_busy
//
// This is a wire, designed to be true is we are ever busy above.
// originally, this was going to be true if we were ever not in the
// idle state.  The logic has since become more complex, hence we have
// a register dedicated to this and just copy out that registers value.
assign	o_busy = (r_busy);


// lcl_data
//
// This is our working copy of the i_data register which we use
// when transmitting.  It is only of interest during transmit, and is
// allowed to be whatever at any other time.  Hence, if r_busy isn't
// true, we can always set it.  On the one clock where r_busy isn't
// true and i_wr is, we set it and r_busy is true thereafter.
// Then, on any zero_baud_counter (i.e. change between baud intervals)
// we simple logically shift the register right to grab the next bit.
initial	lcl_data = 8'hff;
always @(posedge i_clk)
	if ((i_wr)&&(!r_busy))
		lcl_data <= i_data;
	else if (zero_baud_counter)
		lcl_data <= { 1'b1, lcl_data[7:1] };

// o_uart_tx
//
// This is the final result/output desired of this core.  It's all
// centered about o_uart_tx.  This is what finally needs to follow
// the UART protocol.
//
initial	o_uart_tx = 1'b1;
always @(posedge i_clk)
	if ((i_wr)&&(!r_busy))
		o_uart_tx <= 1'b0;	// Set the start bit on writes
	else if (zero_baud_counter)	// Set the data bit.
		o_uart_tx <= lcl_data[0];


// All of the above logic is driven by the baud counter.  Bits must last
// CLOCKS_PER_BAUD in length, and this baud counter is what we use to
// make certain of that.
//
// The basic logic is this: at the beginning of a bit interval, start
// the baud counter and set it to count CLOCKS_PER_BAUD.  When it gets
// to zero, restart it.
//
// However, comparing a 28'bit number to zero can be rather complex--
// especially if we wish to do anything else on that same clock.  For
// that reason, we create "zero_baud_counter".  zero_baud_counter is
// nothing more than a flag that is true anytime baud_counter is zero.
// It's true when the logic (above) needs to step to the next bit.
// Simple enough?
//
// I wish we could stop there, but there are some other (ugly)
// conditions to deal with that offer exceptions to this basic logic.
//
// 1. When the user has commanded a BREAK across the line, we need to
// wait several baud intervals following the break before we start
// transmitting, to give any receiver a chance to recognize that we are
// out of the break condition, and to know that the next bit will be
// a stop bit.
//
// 2. A reset is similar to a break condition--on both we wait several
// baud intervals before allowing a start bit.
//
// 3. In the idle state, we stop our counter--so that upon a request
// to transmit when idle we can start transmitting immediately, rather
// than waiting for the end of the next (fictitious and arbitrary) baud
// interval.
//
// When (i_wr)&&(!r_busy)&&(state == `TXUL_IDLE) then we're not only in
// the idle state, but we also just accepted a command to start writing
// the next word.  At this point, the baud counter needs to be reset
// to the number of CLOCKS_PER_BAUD, and zero_baud_counter set to zero.
//
// The logic is a bit twisted here, in that it will only check for the
// above condition when zero_baud_counter is false--so as to make
// certain the STOP bit is complete.
initial	zero_baud_counter = 1'b1;
initial	baud_counter = 0;
always @(posedge i_clk)
begin
	zero_baud_counter <= (baud_counter == 24'h01);
	if (state == `TXUL_IDLE)
	begin
		baud_counter <= 24'h0;
		zero_baud_counter <= 1'b1;
		if ((i_wr)&&(!r_busy))
		begin
			baud_counter <= CLOCKS_PER_BAUD - 24'h01;
			zero_baud_counter <= 1'b0;
		end
	end else if ((zero_baud_counter)&&(state == 4'h9))
	begin
		baud_counter <= 0;
		zero_baud_counter <= 1'b1;
	end else if (!zero_baud_counter)
		baud_counter <= baud_counter - 24'h01;
	else
		baud_counter <= CLOCKS_PER_BAUD - 24'h01;
end

//
//
// FORMAL METHODS
//
//
//
`ifdef	FORMAL

`ifdef	TXUARTLITE
`define	ASSUME	assume
`else
`define	ASSUME	assert
`endif

// Setup

reg	f_past_valid, f_last_clk;

generate if (F_OPT_CLK2FFLOGIC)
begin

	always @($global_clock)
	begin
		restrict(i_clk == !f_last_clk);
		f_last_clk <= i_clk;
		if (!$rose(i_clk))
		begin
			`ASSUME($stable(i_wr));
			`ASSUME($stable(i_data));
		end
	end

end endgenerate

initial	f_past_valid = 1'b0;
always @(posedge i_clk)
	f_past_valid <= 1'b1;

initial	`ASSUME(!i_wr);
always @(posedge i_clk)
	if ((f_past_valid)&&($past(i_wr))&&($past(o_busy)))
	begin
		`ASSUME(i_wr   == $past(i_wr));
		`ASSUME(i_data == $past(i_data));
	end

// Check the baud counter
always @(posedge i_clk)
	assert(zero_baud_counter == (baud_counter == 0));

always @(posedge i_clk)
	if ((f_past_valid)&&($past(baud_counter != 0))&&($past(state != `TXUL_IDLE)))
		assert(baud_counter == $past(baud_counter - 1'b1));

always @(posedge i_clk)
	if ((f_past_valid)&&(!$past(zero_baud_counter))&&($past(state != `TXUL_IDLE)))
		assert($stable(o_uart_tx));

reg	[(TB-1):0]	f_baud_count;
initial	f_baud_count = 1'b0;
always @(posedge i_clk)
	if (zero_baud_counter)
		f_baud_count <= 0;
	else
		f_baud_count <= f_baud_count + 1'b1;

always @(posedge i_clk)
	assert(f_baud_count < CLOCKS_PER_BAUD);

always @(posedge i_clk)
	if (baud_counter != 0)
		assert(o_busy);

reg	[9:0]	f_txbits;
initial	f_txbits = 0;
always @(posedge i_clk)
	if (zero_baud_counter)
		f_txbits <= { o_uart_tx, f_txbits[9:1] };

always @(posedge i_clk)
if ((f_past_valid)&&(!$past(zero_baud_counter))
		&&(!$past(state==`TXUL_IDLE)))
	assert(state == $past(state));

reg	[3:0]	f_bitcount;
initial	f_bitcount = 0;
always @(posedge i_clk)
	if ((!f_past_valid)||(!$past(f_past_valid)))
		f_bitcount <= 0;
	else if ((state == `TXUL_IDLE)&&(zero_baud_counter))
		f_bitcount <= 0;
	else if (zero_baud_counter)
		f_bitcount <= f_bitcount + 1'b1;

always @(posedge i_clk)
	assert(f_bitcount <= 4'ha);

reg	[7:0]	f_request_tx_data;
always @(posedge i_clk)
	if ((i_wr)&&(!o_busy))
		f_request_tx_data <= i_data;

wire	[3:0]	subcount;
assign	subcount = 10-f_bitcount;
always @(posedge i_clk)
	if (f_bitcount > 0)
		assert(!f_txbits[subcount]);

always @(posedge i_clk)
	if (f_bitcount == 4'ha)
	begin
		assert(f_txbits[8:1] == f_request_tx_data);
		assert( f_txbits[9]);
	end

always @(posedge i_clk)
	assert((state <= `TXUL_STOP + 1'b1)||(state == `TXUL_IDLE));

always @(posedge i_clk)
if ((f_past_valid)&&($past(f_past_valid))&&($past(o_busy)))
	cover(!o_busy);

`endif	// FORMAL
`ifdef	VERIFIC_SVA
reg	[7:0]	fsv_data;

//
// Grab a copy of the data any time we are sent a new byte to transmit
// We'll use this in a moment to compare the item transmitted against
// what is supposed to be transmitted
//
always @(posedge i_clk)
	if ((i_wr)&&(!o_busy))
		fsv_data <= i_data;

//
// One baud interval
//
// 1. The UART output is constant at DAT
// 2. The internal state remains constant at ST
// 3. CKS = the number of clocks per bit.
//
// Everything stays constant during the CKS clocks with the exception
// of (zero_baud_counter), which is *only* raised on the last clock
// interval
sequence	BAUD_INTERVAL(CKS, DAT, SR, ST);
	((o_uart_tx == DAT)&&(state == ST)
		&&(lcl_data == SR)
		&&(!zero_baud_counter))[*(CKS-1)]
	##1 (o_uart_tx == DAT)&&(state == ST)
		&&(lcl_data == SR)
		&&(zero_baud_counter);
endsequence

//
// One byte transmitted
//
// DATA = the byte that is sent
// CKS  = the number of clocks per bit
//
sequence	SEND(CKS, DATA);
	BAUD_INTERVAL(CKS, 1'b0, DATA, 4'h0)
	##1 BAUD_INTERVAL(CKS, DATA[0], {{(1){1'b1}},DATA[7:1]}, 4'h1)
	##1 BAUD_INTERVAL(CKS, DATA[1], {{(2){1'b1}},DATA[7:2]}, 4'h2)
	##1 BAUD_INTERVAL(CKS, DATA[2], {{(3){1'b1}},DATA[7:3]}, 4'h3)
	##1 BAUD_INTERVAL(CKS, DATA[3], {{(4){1'b1}},DATA[7:4]}, 4'h4)
	##1 BAUD_INTERVAL(CKS, DATA[4], {{(5){1'b1}},DATA[7:5]}, 4'h5)
	##1 BAUD_INTERVAL(CKS, DATA[5], {{(6){1'b1}},DATA[7:6]}, 4'h6)
	##1 BAUD_INTERVAL(CKS, DATA[6], {{(7){1'b1}},DATA[7:7]}, 4'h7)
	##1 BAUD_INTERVAL(CKS, DATA[7], 8'hff, 4'h8)
	##1 BAUD_INTERVAL(CKS, 1'b1, 8'hff, 4'h9);
endsequence

//
// Transmit one byte
//
// Once the byte is transmitted, make certain we return to
// idle
//
assert property (
	@(posedge i_clk)
	(i_wr)&&(!o_busy)
	|=> ((o_busy) throughout SEND(CLOCKS_PER_BAUD,fsv_data))
	##1 (!o_busy)&&(o_uart_tx)&&(zero_baud_counter));

assume property (
	@(posedge i_clk)
	(i_wr)&&(o_busy) |=>
		(i_wr)&&(o_busy)&&($stable(i_data)));

//
// Make certain that o_busy is true any time zero_baud_counter is
// non-zero
//
always @(*)
	assert((o_busy)||(zero_baud_counter) );

// If and only if zero_baud_counter is true, baud_counter must be zero
// Insist on that relationship here.
always @(*)
	assert(zero_baud_counter == (baud_counter == 0));

// To make certain baud_counter stays below CLOCKS_PER_BAUD
always @(*)
	assert(baud_counter < CLOCKS_PER_BAUD);

//
// Insist that we are only ever in a valid state
always @(*)
	assert((state <= `TXUL_STOP+1'b1)||(state == `TXUL_IDLE));

`endif // Verific SVA
endmodule